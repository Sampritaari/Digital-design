magic
tech sky130A
magscale 1 2
timestamp 1755980430
<< viali >>
rect 4721 10217 4755 10251
rect 6745 10217 6779 10251
rect 2513 10149 2547 10183
rect 1501 10013 1535 10047
rect 2973 10013 3007 10047
rect 6653 10013 6687 10047
rect 8033 10013 8067 10047
rect 8309 10013 8343 10047
rect 8585 10013 8619 10047
rect 1685 9945 1719 9979
rect 2697 9945 2731 9979
rect 4997 9945 5031 9979
rect 7481 9945 7515 9979
rect 7665 9945 7699 9979
rect 3065 9877 3099 9911
rect 7941 9877 7975 9911
rect 8401 9877 8435 9911
rect 8769 9877 8803 9911
rect 4813 9673 4847 9707
rect 8585 9673 8619 9707
rect 2973 9605 3007 9639
rect 3617 9605 3651 9639
rect 3801 9605 3835 9639
rect 3985 9605 4019 9639
rect 4721 9605 4755 9639
rect 6745 9605 6779 9639
rect 8677 9605 8711 9639
rect 1409 9537 1443 9571
rect 2329 9537 2363 9571
rect 2421 9537 2455 9571
rect 2605 9537 2639 9571
rect 2697 9537 2731 9571
rect 2789 9537 2823 9571
rect 3065 9537 3099 9571
rect 3157 9537 3191 9571
rect 3893 9537 3927 9571
rect 4169 9537 4203 9571
rect 4445 9537 4479 9571
rect 4997 9537 5031 9571
rect 5089 9537 5123 9571
rect 5181 9537 5215 9571
rect 5365 9537 5399 9571
rect 5457 9537 5491 9571
rect 5549 9537 5583 9571
rect 5734 9537 5768 9571
rect 5825 9537 5859 9571
rect 6101 9537 6135 9571
rect 6653 9537 6687 9571
rect 6929 9537 6963 9571
rect 7021 9537 7055 9571
rect 7297 9537 7331 9571
rect 7389 9537 7423 9571
rect 7849 9537 7883 9571
rect 1685 9469 1719 9503
rect 4353 9469 4387 9503
rect 4721 9469 4755 9503
rect 7573 9469 7607 9503
rect 7757 9469 7791 9503
rect 7941 9469 7975 9503
rect 8033 9469 8067 9503
rect 8217 9469 8251 9503
rect 3617 9401 3651 9435
rect 6929 9401 6963 9435
rect 2605 9333 2639 9367
rect 3341 9333 3375 9367
rect 4537 9333 4571 9367
rect 6009 9333 6043 9367
rect 7113 9333 7147 9367
rect 2881 9129 2915 9163
rect 4353 9129 4387 9163
rect 5825 9129 5859 9163
rect 2421 9061 2455 9095
rect 8309 9061 8343 9095
rect 8033 8993 8067 9027
rect 1409 8925 1443 8959
rect 1685 8925 1719 8959
rect 2329 8925 2363 8959
rect 2605 8925 2639 8959
rect 2697 8925 2731 8959
rect 3801 8925 3835 8959
rect 4169 8925 4203 8959
rect 4261 8925 4295 8959
rect 4445 8925 4479 8959
rect 5549 8925 5583 8959
rect 7941 8925 7975 8959
rect 8769 8925 8803 8959
rect 3985 8857 4019 8891
rect 5825 8857 5859 8891
rect 5641 8789 5675 8823
rect 8585 8789 8619 8823
rect 2237 8585 2271 8619
rect 5273 8585 5307 8619
rect 7113 8585 7147 8619
rect 8309 8585 8343 8619
rect 4169 8517 4203 8551
rect 4261 8517 4295 8551
rect 6745 8517 6779 8551
rect 7665 8517 7699 8551
rect 1869 8449 1903 8483
rect 2973 8449 3007 8483
rect 3985 8449 4019 8483
rect 4353 8449 4387 8483
rect 5181 8449 5215 8483
rect 5365 8449 5399 8483
rect 6929 8449 6963 8483
rect 7205 8449 7239 8483
rect 7481 8449 7515 8483
rect 7757 8449 7791 8483
rect 7849 8449 7883 8483
rect 8677 8449 8711 8483
rect 1777 8381 1811 8415
rect 3249 8381 3283 8415
rect 4537 8313 4571 8347
rect 7297 8313 7331 8347
rect 8953 8313 8987 8347
rect 2789 8245 2823 8279
rect 3157 8245 3191 8279
rect 7941 8245 7975 8279
rect 1961 8041 1995 8075
rect 5089 8041 5123 8075
rect 6929 8041 6963 8075
rect 7481 8041 7515 8075
rect 7573 8041 7607 8075
rect 7757 8041 7791 8075
rect 8033 8041 8067 8075
rect 8401 8041 8435 8075
rect 5641 7973 5675 8007
rect 2697 7905 2731 7939
rect 3617 7905 3651 7939
rect 4537 7905 4571 7939
rect 4997 7905 5031 7939
rect 6009 7905 6043 7939
rect 2145 7837 2179 7871
rect 2421 7837 2455 7871
rect 2973 7837 3007 7871
rect 4629 7837 4663 7871
rect 5273 7837 5307 7871
rect 5549 7837 5583 7871
rect 5825 7837 5859 7871
rect 6285 7837 6319 7871
rect 6653 7837 6687 7871
rect 6745 7837 6779 7871
rect 7095 7837 7129 7871
rect 7205 7837 7239 7871
rect 7297 7837 7331 7871
rect 8493 7837 8527 7871
rect 2329 7769 2363 7803
rect 7725 7769 7759 7803
rect 7941 7769 7975 7803
rect 5457 7701 5491 7735
rect 5273 7497 5307 7531
rect 8861 7497 8895 7531
rect 1777 7361 1811 7395
rect 2697 7361 2731 7395
rect 2881 7361 2915 7395
rect 3157 7361 3191 7395
rect 5457 7361 5491 7395
rect 5549 7361 5583 7395
rect 8677 7361 8711 7395
rect 2973 7293 3007 7327
rect 5273 7293 5307 7327
rect 8401 7293 8435 7327
rect 2789 7225 2823 7259
rect 8493 7225 8527 7259
rect 1501 7157 1535 7191
rect 2421 7157 2455 7191
rect 7941 6885 7975 6919
rect 1777 6817 1811 6851
rect 2053 6817 2087 6851
rect 3801 6817 3835 6851
rect 1685 6749 1719 6783
rect 3985 6749 4019 6783
rect 4353 6749 4387 6783
rect 7297 6749 7331 6783
rect 7665 6749 7699 6783
rect 7941 6749 7975 6783
rect 8401 6749 8435 6783
rect 3893 6681 3927 6715
rect 4629 6681 4663 6715
rect 8125 6681 8159 6715
rect 7481 6613 7515 6647
rect 8223 6613 8257 6647
rect 8309 6613 8343 6647
rect 2237 6409 2271 6443
rect 6009 6409 6043 6443
rect 7113 6409 7147 6443
rect 8677 6409 8711 6443
rect 2605 6341 2639 6375
rect 6754 6341 6788 6375
rect 2148 6295 2182 6329
rect 2421 6273 2455 6307
rect 3617 6273 3651 6307
rect 3801 6273 3835 6307
rect 3893 6273 3927 6307
rect 4077 6273 4111 6307
rect 4445 6273 4479 6307
rect 4629 6273 4663 6307
rect 4721 6273 4755 6307
rect 4813 6273 4847 6307
rect 6193 6273 6227 6307
rect 6377 6273 6411 6307
rect 7389 6273 7423 6307
rect 7665 6273 7699 6307
rect 7941 6273 7975 6307
rect 8034 6273 8068 6307
rect 8217 6273 8251 6307
rect 8309 6273 8343 6307
rect 8406 6273 8440 6307
rect 8953 6273 8987 6307
rect 4353 6205 4387 6239
rect 8677 6205 8711 6239
rect 8585 6137 8619 6171
rect 3433 6069 3467 6103
rect 4261 6069 4295 6103
rect 5089 6069 5123 6103
rect 6745 6069 6779 6103
rect 6929 6069 6963 6103
rect 7573 6069 7607 6103
rect 8861 6069 8895 6103
rect 2789 5865 2823 5899
rect 4997 5865 5031 5899
rect 7113 5865 7147 5899
rect 7297 5865 7331 5899
rect 7849 5865 7883 5899
rect 8217 5865 8251 5899
rect 8677 5865 8711 5899
rect 2237 5797 2271 5831
rect 1961 5729 1995 5763
rect 2421 5729 2455 5763
rect 3985 5729 4019 5763
rect 4261 5729 4295 5763
rect 4813 5729 4847 5763
rect 1777 5661 1811 5695
rect 1869 5661 1903 5695
rect 2053 5661 2087 5695
rect 2513 5661 2547 5695
rect 4077 5661 4111 5695
rect 4169 5661 4203 5695
rect 5089 5661 5123 5695
rect 7389 5661 7423 5695
rect 7665 5661 7699 5695
rect 7757 5661 7791 5695
rect 8493 5661 8527 5695
rect 4445 5525 4479 5559
rect 4813 5525 4847 5559
rect 1777 5321 1811 5355
rect 8033 5321 8067 5355
rect 1685 5253 1719 5287
rect 2697 5253 2731 5287
rect 1409 5185 1443 5219
rect 1501 5185 1535 5219
rect 1961 5185 1995 5219
rect 2053 5185 2087 5219
rect 2329 5185 2363 5219
rect 2881 5185 2915 5219
rect 4629 5185 4663 5219
rect 5089 5185 5123 5219
rect 5273 5185 5307 5219
rect 5365 5185 5399 5219
rect 5457 5185 5491 5219
rect 7665 5185 7699 5219
rect 8769 5185 8803 5219
rect 4537 5117 4571 5151
rect 7573 5117 7607 5151
rect 7757 5117 7791 5151
rect 7849 5117 7883 5151
rect 9045 5117 9079 5151
rect 1685 5049 1719 5083
rect 2237 5049 2271 5083
rect 3065 4981 3099 5015
rect 4905 4981 4939 5015
rect 5733 4981 5767 5015
rect 2605 4777 2639 4811
rect 5457 4777 5491 4811
rect 7205 4777 7239 4811
rect 7573 4777 7607 4811
rect 1685 4709 1719 4743
rect 6745 4709 6779 4743
rect 8217 4709 8251 4743
rect 4813 4641 4847 4675
rect 5641 4641 5675 4675
rect 6929 4641 6963 4675
rect 7297 4641 7331 4675
rect 1501 4573 1535 4607
rect 2513 4573 2547 4607
rect 3801 4573 3835 4607
rect 3985 4573 4019 4607
rect 4077 4573 4111 4607
rect 4261 4573 4295 4607
rect 4997 4573 5031 4607
rect 5273 4573 5307 4607
rect 5733 4573 5767 4607
rect 7205 4573 7239 4607
rect 7941 4573 7975 4607
rect 8125 4573 8159 4607
rect 6469 4505 6503 4539
rect 3801 4437 3835 4471
rect 4261 4437 4295 4471
rect 5181 4437 5215 4471
rect 1685 4097 1719 4131
rect 1869 4097 1903 4131
rect 2053 4097 2087 4131
rect 2145 4097 2179 4131
rect 2881 4097 2915 4131
rect 3065 4097 3099 4131
rect 3341 4097 3375 4131
rect 3525 4097 3559 4131
rect 3893 4097 3927 4131
rect 7021 4097 7055 4131
rect 3617 4029 3651 4063
rect 3709 4029 3743 4063
rect 4077 4029 4111 4063
rect 7113 4029 7147 4063
rect 7297 4029 7331 4063
rect 3157 3961 3191 3995
rect 7205 3961 7239 3995
rect 2973 3893 3007 3927
rect 1593 3689 1627 3723
rect 1777 3689 1811 3723
rect 3525 3689 3559 3723
rect 5089 3689 5123 3723
rect 4353 3621 4387 3655
rect 8493 3621 8527 3655
rect 1961 3553 1995 3587
rect 2145 3553 2179 3587
rect 5457 3553 5491 3587
rect 7389 3553 7423 3587
rect 7665 3553 7699 3587
rect 2053 3485 2087 3519
rect 2237 3485 2271 3519
rect 4353 3485 4387 3519
rect 4629 3485 4663 3519
rect 5273 3485 5307 3519
rect 5365 3485 5399 3519
rect 5549 3485 5583 3519
rect 7757 3485 7791 3519
rect 8677 3485 8711 3519
rect 1501 3417 1535 3451
rect 3157 3417 3191 3451
rect 3341 3417 3375 3451
rect 4537 3349 4571 3383
rect 1777 3145 1811 3179
rect 2513 3145 2547 3179
rect 3433 3145 3467 3179
rect 5917 3145 5951 3179
rect 7205 3145 7239 3179
rect 7849 3145 7883 3179
rect 8125 3145 8159 3179
rect 1593 3077 1627 3111
rect 3617 3077 3651 3111
rect 5273 3077 5307 3111
rect 1869 3009 1903 3043
rect 1961 3009 1995 3043
rect 2237 3009 2271 3043
rect 2329 3009 2363 3043
rect 2789 3009 2823 3043
rect 3249 3009 3283 3043
rect 3433 3009 3467 3043
rect 3525 3009 3559 3043
rect 4261 3009 4295 3043
rect 4813 3009 4847 3043
rect 4905 3009 4939 3043
rect 5089 3009 5123 3043
rect 5365 3009 5399 3043
rect 5641 3009 5675 3043
rect 5733 3009 5767 3043
rect 6837 3009 6871 3043
rect 7297 3009 7331 3043
rect 7573 3009 7607 3043
rect 7665 3009 7699 3043
rect 7941 3009 7975 3043
rect 8769 3009 8803 3043
rect 8953 3009 8987 3043
rect 2881 2941 2915 2975
rect 3157 2941 3191 2975
rect 4353 2941 4387 2975
rect 6929 2941 6963 2975
rect 1593 2873 1627 2907
rect 2053 2873 2087 2907
rect 4997 2873 5031 2907
rect 5457 2873 5491 2907
rect 4537 2805 4571 2839
rect 7389 2805 7423 2839
rect 2513 2601 2547 2635
rect 5733 2601 5767 2635
rect 6009 2601 6043 2635
rect 7389 2601 7423 2635
rect 8585 2601 8619 2635
rect 1685 2533 1719 2567
rect 4077 2533 4111 2567
rect 8033 2533 8067 2567
rect 2973 2465 3007 2499
rect 7757 2465 7791 2499
rect 7849 2465 7883 2499
rect 2329 2397 2363 2431
rect 2697 2397 2731 2431
rect 5457 2397 5491 2431
rect 5549 2397 5583 2431
rect 6653 2397 6687 2431
rect 7573 2397 7607 2431
rect 7665 2397 7699 2431
rect 8217 2397 8251 2431
rect 8309 2397 8343 2431
rect 1501 2329 1535 2363
rect 3893 2329 3927 2363
rect 5733 2329 5767 2363
rect 5917 2329 5951 2363
rect 8033 2329 8067 2363
rect 8677 2329 8711 2363
rect 6929 2261 6963 2295
<< metal1 >>
rect 1104 10362 9384 10384
rect 1104 10310 1985 10362
rect 2037 10310 2049 10362
rect 2101 10310 2113 10362
rect 2165 10310 2177 10362
rect 2229 10310 2241 10362
rect 2293 10310 4055 10362
rect 4107 10310 4119 10362
rect 4171 10310 4183 10362
rect 4235 10310 4247 10362
rect 4299 10310 4311 10362
rect 4363 10310 6125 10362
rect 6177 10310 6189 10362
rect 6241 10310 6253 10362
rect 6305 10310 6317 10362
rect 6369 10310 6381 10362
rect 6433 10310 8195 10362
rect 8247 10310 8259 10362
rect 8311 10310 8323 10362
rect 8375 10310 8387 10362
rect 8439 10310 8451 10362
rect 8503 10310 9384 10362
rect 1104 10288 9384 10310
rect 4614 10208 4620 10260
rect 4672 10248 4678 10260
rect 4709 10251 4767 10257
rect 4709 10248 4721 10251
rect 4672 10220 4721 10248
rect 4672 10208 4678 10220
rect 4709 10217 4721 10220
rect 4755 10217 4767 10251
rect 4709 10211 4767 10217
rect 6730 10208 6736 10260
rect 6788 10208 6794 10260
rect 2501 10183 2559 10189
rect 2501 10149 2513 10183
rect 2547 10180 2559 10183
rect 2774 10180 2780 10192
rect 2547 10152 2780 10180
rect 2547 10149 2559 10152
rect 2501 10143 2559 10149
rect 2774 10140 2780 10152
rect 2832 10140 2838 10192
rect 1302 10004 1308 10056
rect 1360 10044 1366 10056
rect 1489 10047 1547 10053
rect 1489 10044 1501 10047
rect 1360 10016 1501 10044
rect 1360 10004 1366 10016
rect 1489 10013 1501 10016
rect 1535 10013 1547 10047
rect 1489 10007 1547 10013
rect 2590 10004 2596 10056
rect 2648 10044 2654 10056
rect 2961 10047 3019 10053
rect 2961 10044 2973 10047
rect 2648 10016 2973 10044
rect 2648 10004 2654 10016
rect 2961 10013 2973 10016
rect 3007 10013 3019 10047
rect 2961 10007 3019 10013
rect 4154 10004 4160 10056
rect 4212 10044 4218 10056
rect 6641 10047 6699 10053
rect 6641 10044 6653 10047
rect 4212 10016 6653 10044
rect 4212 10004 4218 10016
rect 6641 10013 6653 10016
rect 6687 10013 6699 10047
rect 6641 10007 6699 10013
rect 7742 10004 7748 10056
rect 7800 10044 7806 10056
rect 8021 10047 8079 10053
rect 8021 10044 8033 10047
rect 7800 10016 8033 10044
rect 7800 10004 7806 10016
rect 8021 10013 8033 10016
rect 8067 10013 8079 10047
rect 8021 10007 8079 10013
rect 8297 10047 8355 10053
rect 8297 10013 8309 10047
rect 8343 10044 8355 10047
rect 8478 10044 8484 10056
rect 8343 10016 8484 10044
rect 8343 10013 8355 10016
rect 8297 10007 8355 10013
rect 8478 10004 8484 10016
rect 8536 10004 8542 10056
rect 8573 10047 8631 10053
rect 8573 10013 8585 10047
rect 8619 10044 8631 10047
rect 8662 10044 8668 10056
rect 8619 10016 8668 10044
rect 8619 10013 8631 10016
rect 8573 10007 8631 10013
rect 8662 10004 8668 10016
rect 8720 10004 8726 10056
rect 9674 10004 9680 10056
rect 9732 10004 9738 10056
rect 1670 9936 1676 9988
rect 1728 9936 1734 9988
rect 2498 9936 2504 9988
rect 2556 9976 2562 9988
rect 2685 9979 2743 9985
rect 2685 9976 2697 9979
rect 2556 9948 2697 9976
rect 2556 9936 2562 9948
rect 2685 9945 2697 9948
rect 2731 9945 2743 9979
rect 2685 9939 2743 9945
rect 4985 9979 5043 9985
rect 4985 9945 4997 9979
rect 5031 9976 5043 9979
rect 5074 9976 5080 9988
rect 5031 9948 5080 9976
rect 5031 9945 5043 9948
rect 4985 9939 5043 9945
rect 5074 9936 5080 9948
rect 5132 9936 5138 9988
rect 7282 9936 7288 9988
rect 7340 9976 7346 9988
rect 7469 9979 7527 9985
rect 7469 9976 7481 9979
rect 7340 9948 7481 9976
rect 7340 9936 7346 9948
rect 7469 9945 7481 9948
rect 7515 9945 7527 9979
rect 7469 9939 7527 9945
rect 7653 9979 7711 9985
rect 7653 9945 7665 9979
rect 7699 9976 7711 9979
rect 9692 9976 9720 10004
rect 7699 9948 9720 9976
rect 7699 9945 7711 9948
rect 7653 9939 7711 9945
rect 3053 9911 3111 9917
rect 3053 9877 3065 9911
rect 3099 9908 3111 9911
rect 6638 9908 6644 9920
rect 3099 9880 6644 9908
rect 3099 9877 3111 9880
rect 3053 9871 3111 9877
rect 6638 9868 6644 9880
rect 6696 9868 6702 9920
rect 7926 9868 7932 9920
rect 7984 9868 7990 9920
rect 8386 9868 8392 9920
rect 8444 9868 8450 9920
rect 8754 9868 8760 9920
rect 8812 9868 8818 9920
rect 1104 9818 9384 9840
rect 1104 9766 2645 9818
rect 2697 9766 2709 9818
rect 2761 9766 2773 9818
rect 2825 9766 2837 9818
rect 2889 9766 2901 9818
rect 2953 9766 4715 9818
rect 4767 9766 4779 9818
rect 4831 9766 4843 9818
rect 4895 9766 4907 9818
rect 4959 9766 4971 9818
rect 5023 9766 6785 9818
rect 6837 9766 6849 9818
rect 6901 9766 6913 9818
rect 6965 9766 6977 9818
rect 7029 9766 7041 9818
rect 7093 9766 8855 9818
rect 8907 9766 8919 9818
rect 8971 9766 8983 9818
rect 9035 9766 9047 9818
rect 9099 9766 9111 9818
rect 9163 9766 9384 9818
rect 1104 9744 9384 9766
rect 4801 9707 4859 9713
rect 3712 9676 4568 9704
rect 2961 9639 3019 9645
rect 2961 9636 2973 9639
rect 2424 9608 2973 9636
rect 1394 9528 1400 9580
rect 1452 9528 1458 9580
rect 2314 9528 2320 9580
rect 2372 9528 2378 9580
rect 2424 9577 2452 9608
rect 2961 9605 2973 9608
rect 3007 9636 3019 9639
rect 3605 9639 3663 9645
rect 3007 9608 3556 9636
rect 3007 9605 3019 9608
rect 2961 9599 3019 9605
rect 2409 9571 2467 9577
rect 2409 9537 2421 9571
rect 2455 9537 2467 9571
rect 2409 9531 2467 9537
rect 2593 9571 2651 9577
rect 2593 9537 2605 9571
rect 2639 9537 2651 9571
rect 2593 9531 2651 9537
rect 1670 9460 1676 9512
rect 1728 9460 1734 9512
rect 2424 9500 2452 9531
rect 1780 9472 2452 9500
rect 1780 9444 1808 9472
rect 1762 9392 1768 9444
rect 1820 9392 1826 9444
rect 2608 9432 2636 9531
rect 2682 9528 2688 9580
rect 2740 9528 2746 9580
rect 2777 9571 2835 9577
rect 2777 9537 2789 9571
rect 2823 9537 2835 9571
rect 2777 9531 2835 9537
rect 2792 9500 2820 9531
rect 3050 9528 3056 9580
rect 3108 9528 3114 9580
rect 3145 9571 3203 9577
rect 3145 9537 3157 9571
rect 3191 9568 3203 9571
rect 3234 9568 3240 9580
rect 3191 9540 3240 9568
rect 3191 9537 3203 9540
rect 3145 9531 3203 9537
rect 3234 9528 3240 9540
rect 3292 9528 3298 9580
rect 3528 9568 3556 9608
rect 3605 9605 3617 9639
rect 3651 9636 3663 9639
rect 3712 9636 3740 9676
rect 3651 9608 3740 9636
rect 3789 9639 3847 9645
rect 3651 9605 3663 9608
rect 3605 9599 3663 9605
rect 3789 9605 3801 9639
rect 3835 9636 3847 9639
rect 3973 9639 4031 9645
rect 3973 9636 3985 9639
rect 3835 9608 3985 9636
rect 3835 9605 3847 9608
rect 3789 9599 3847 9605
rect 3973 9605 3985 9608
rect 4019 9636 4031 9639
rect 4540 9636 4568 9676
rect 4801 9673 4813 9707
rect 4847 9704 4859 9707
rect 5074 9704 5080 9716
rect 4847 9676 5080 9704
rect 4847 9673 4859 9676
rect 4801 9667 4859 9673
rect 5074 9664 5080 9676
rect 5132 9664 5138 9716
rect 8386 9704 8392 9716
rect 5184 9676 8392 9704
rect 4709 9639 4767 9645
rect 4709 9636 4721 9639
rect 4019 9608 4476 9636
rect 4540 9608 4721 9636
rect 4019 9605 4031 9608
rect 3973 9599 4031 9605
rect 3881 9571 3939 9577
rect 3528 9540 3832 9568
rect 3804 9512 3832 9540
rect 3881 9537 3893 9571
rect 3927 9568 3939 9571
rect 4062 9568 4068 9580
rect 3927 9540 4068 9568
rect 3927 9537 3939 9540
rect 3881 9531 3939 9537
rect 4062 9528 4068 9540
rect 4120 9528 4126 9580
rect 4157 9571 4215 9577
rect 4157 9537 4169 9571
rect 4203 9568 4215 9571
rect 4246 9568 4252 9580
rect 4203 9540 4252 9568
rect 4203 9537 4215 9540
rect 4157 9531 4215 9537
rect 4246 9528 4252 9540
rect 4304 9528 4310 9580
rect 4448 9577 4476 9608
rect 4709 9605 4721 9608
rect 4755 9605 4767 9639
rect 5184 9636 5212 9676
rect 8386 9664 8392 9676
rect 8444 9664 8450 9716
rect 8573 9707 8631 9713
rect 8573 9673 8585 9707
rect 8619 9704 8631 9707
rect 9398 9704 9404 9716
rect 8619 9676 9404 9704
rect 8619 9673 8631 9676
rect 8573 9667 8631 9673
rect 9398 9664 9404 9676
rect 9456 9664 9462 9716
rect 6733 9639 6791 9645
rect 4709 9599 4767 9605
rect 4908 9608 5212 9636
rect 5276 9608 6132 9636
rect 4433 9571 4491 9577
rect 4433 9537 4445 9571
rect 4479 9537 4491 9571
rect 4433 9531 4491 9537
rect 4908 9512 4936 9608
rect 4982 9528 4988 9580
rect 5040 9528 5046 9580
rect 5077 9571 5135 9577
rect 5077 9537 5089 9571
rect 5123 9537 5135 9571
rect 5077 9531 5135 9537
rect 2792 9472 3648 9500
rect 3620 9441 3648 9472
rect 3786 9460 3792 9512
rect 3844 9460 3850 9512
rect 3970 9460 3976 9512
rect 4028 9500 4034 9512
rect 4341 9503 4399 9509
rect 4028 9472 4292 9500
rect 4028 9460 4034 9472
rect 3605 9435 3663 9441
rect 2240 9404 2728 9432
rect 1394 9324 1400 9376
rect 1452 9364 1458 9376
rect 2240 9364 2268 9404
rect 1452 9336 2268 9364
rect 1452 9324 1458 9336
rect 2590 9324 2596 9376
rect 2648 9324 2654 9376
rect 2700 9364 2728 9404
rect 3605 9401 3617 9435
rect 3651 9401 3663 9435
rect 4154 9432 4160 9444
rect 3605 9395 3663 9401
rect 3804 9404 4160 9432
rect 3234 9364 3240 9376
rect 2700 9336 3240 9364
rect 3234 9324 3240 9336
rect 3292 9324 3298 9376
rect 3329 9367 3387 9373
rect 3329 9333 3341 9367
rect 3375 9364 3387 9367
rect 3804 9364 3832 9404
rect 4154 9392 4160 9404
rect 4212 9392 4218 9444
rect 4264 9432 4292 9472
rect 4341 9469 4353 9503
rect 4387 9500 4399 9503
rect 4614 9500 4620 9512
rect 4387 9472 4620 9500
rect 4387 9469 4399 9472
rect 4341 9463 4399 9469
rect 4614 9460 4620 9472
rect 4672 9460 4678 9512
rect 4709 9503 4767 9509
rect 4709 9469 4721 9503
rect 4755 9500 4767 9503
rect 4890 9500 4896 9512
rect 4755 9472 4896 9500
rect 4755 9469 4767 9472
rect 4709 9463 4767 9469
rect 4890 9460 4896 9472
rect 4948 9460 4954 9512
rect 5092 9500 5120 9531
rect 5166 9528 5172 9580
rect 5224 9568 5230 9580
rect 5276 9568 5304 9608
rect 5224 9540 5304 9568
rect 5224 9528 5230 9540
rect 5350 9528 5356 9580
rect 5408 9528 5414 9580
rect 5445 9571 5503 9577
rect 5445 9537 5457 9571
rect 5491 9568 5503 9571
rect 5537 9571 5595 9577
rect 5537 9568 5549 9571
rect 5491 9540 5549 9568
rect 5491 9537 5503 9540
rect 5445 9531 5503 9537
rect 5537 9537 5549 9540
rect 5583 9537 5595 9571
rect 5718 9568 5724 9580
rect 5537 9531 5595 9537
rect 5644 9540 5724 9568
rect 5258 9500 5264 9512
rect 5092 9472 5264 9500
rect 5258 9460 5264 9472
rect 5316 9460 5322 9512
rect 5644 9432 5672 9540
rect 5718 9528 5724 9540
rect 5776 9528 5782 9580
rect 6104 9577 6132 9608
rect 6733 9605 6745 9639
rect 6779 9636 6791 9639
rect 8665 9639 8723 9645
rect 6779 9608 7880 9636
rect 6779 9605 6791 9608
rect 6733 9599 6791 9605
rect 5813 9571 5871 9577
rect 5813 9537 5825 9571
rect 5859 9537 5871 9571
rect 5813 9531 5871 9537
rect 6089 9571 6147 9577
rect 6089 9537 6101 9571
rect 6135 9537 6147 9571
rect 6089 9531 6147 9537
rect 6641 9571 6699 9577
rect 6641 9537 6653 9571
rect 6687 9537 6699 9571
rect 6641 9531 6699 9537
rect 4264 9404 5672 9432
rect 5828 9376 5856 9531
rect 6656 9432 6684 9531
rect 6914 9528 6920 9580
rect 6972 9528 6978 9580
rect 7024 9577 7052 9608
rect 7009 9571 7067 9577
rect 7009 9537 7021 9571
rect 7055 9537 7067 9571
rect 7009 9531 7067 9537
rect 7285 9571 7343 9577
rect 7285 9537 7297 9571
rect 7331 9537 7343 9571
rect 7285 9531 7343 9537
rect 7300 9500 7328 9531
rect 7374 9528 7380 9580
rect 7432 9528 7438 9580
rect 7852 9577 7880 9608
rect 8665 9605 8677 9639
rect 8711 9636 8723 9639
rect 8754 9636 8760 9648
rect 8711 9608 8760 9636
rect 8711 9605 8723 9608
rect 8665 9599 8723 9605
rect 8754 9596 8760 9608
rect 8812 9596 8818 9648
rect 7837 9571 7895 9577
rect 7837 9537 7849 9571
rect 7883 9568 7895 9571
rect 7883 9540 8156 9568
rect 7883 9537 7895 9540
rect 7837 9531 7895 9537
rect 8128 9512 8156 9540
rect 6932 9472 7328 9500
rect 7561 9503 7619 9509
rect 6932 9441 6960 9472
rect 7561 9469 7573 9503
rect 7607 9500 7619 9503
rect 7745 9503 7803 9509
rect 7745 9500 7757 9503
rect 7607 9472 7757 9500
rect 7607 9469 7619 9472
rect 7561 9463 7619 9469
rect 7745 9469 7757 9472
rect 7791 9469 7803 9503
rect 7745 9463 7803 9469
rect 7926 9460 7932 9512
rect 7984 9460 7990 9512
rect 8021 9503 8079 9509
rect 8021 9469 8033 9503
rect 8067 9469 8079 9503
rect 8021 9463 8079 9469
rect 6917 9435 6975 9441
rect 5920 9404 6868 9432
rect 5920 9376 5948 9404
rect 3375 9336 3832 9364
rect 3375 9333 3387 9336
rect 3329 9327 3387 9333
rect 4062 9324 4068 9376
rect 4120 9364 4126 9376
rect 4525 9367 4583 9373
rect 4525 9364 4537 9367
rect 4120 9336 4537 9364
rect 4120 9324 4126 9336
rect 4525 9333 4537 9336
rect 4571 9364 4583 9367
rect 5074 9364 5080 9376
rect 4571 9336 5080 9364
rect 4571 9333 4583 9336
rect 4525 9327 4583 9333
rect 5074 9324 5080 9336
rect 5132 9324 5138 9376
rect 5810 9324 5816 9376
rect 5868 9324 5874 9376
rect 5902 9324 5908 9376
rect 5960 9324 5966 9376
rect 5994 9324 6000 9376
rect 6052 9324 6058 9376
rect 6840 9364 6868 9404
rect 6917 9401 6929 9435
rect 6963 9401 6975 9435
rect 7944 9432 7972 9460
rect 6917 9395 6975 9401
rect 7116 9404 7972 9432
rect 7116 9373 7144 9404
rect 7101 9367 7159 9373
rect 7101 9364 7113 9367
rect 6840 9336 7113 9364
rect 7101 9333 7113 9336
rect 7147 9333 7159 9367
rect 7101 9327 7159 9333
rect 7742 9324 7748 9376
rect 7800 9364 7806 9376
rect 8036 9364 8064 9463
rect 8110 9460 8116 9512
rect 8168 9460 8174 9512
rect 8205 9503 8263 9509
rect 8205 9469 8217 9503
rect 8251 9500 8263 9503
rect 8662 9500 8668 9512
rect 8251 9472 8668 9500
rect 8251 9469 8263 9472
rect 8205 9463 8263 9469
rect 8662 9460 8668 9472
rect 8720 9460 8726 9512
rect 7800 9336 8064 9364
rect 7800 9324 7806 9336
rect 1104 9274 9384 9296
rect 1104 9222 1985 9274
rect 2037 9222 2049 9274
rect 2101 9222 2113 9274
rect 2165 9222 2177 9274
rect 2229 9222 2241 9274
rect 2293 9222 4055 9274
rect 4107 9222 4119 9274
rect 4171 9222 4183 9274
rect 4235 9222 4247 9274
rect 4299 9222 4311 9274
rect 4363 9222 6125 9274
rect 6177 9222 6189 9274
rect 6241 9222 6253 9274
rect 6305 9222 6317 9274
rect 6369 9222 6381 9274
rect 6433 9222 8195 9274
rect 8247 9222 8259 9274
rect 8311 9222 8323 9274
rect 8375 9222 8387 9274
rect 8439 9222 8451 9274
rect 8503 9222 9384 9274
rect 1104 9200 9384 9222
rect 2590 9120 2596 9172
rect 2648 9120 2654 9172
rect 2682 9120 2688 9172
rect 2740 9160 2746 9172
rect 2869 9163 2927 9169
rect 2869 9160 2881 9163
rect 2740 9132 2881 9160
rect 2740 9120 2746 9132
rect 2869 9129 2881 9132
rect 2915 9129 2927 9163
rect 2869 9123 2927 9129
rect 3234 9120 3240 9172
rect 3292 9160 3298 9172
rect 4341 9163 4399 9169
rect 3292 9132 4108 9160
rect 3292 9120 3298 9132
rect 2409 9095 2467 9101
rect 2409 9061 2421 9095
rect 2455 9061 2467 9095
rect 2409 9055 2467 9061
rect 2424 8968 2452 9055
rect 934 8916 940 8968
rect 992 8956 998 8968
rect 1397 8959 1455 8965
rect 1397 8956 1409 8959
rect 992 8928 1409 8956
rect 992 8916 998 8928
rect 1397 8925 1409 8928
rect 1443 8925 1455 8959
rect 1397 8919 1455 8925
rect 1673 8959 1731 8965
rect 1673 8925 1685 8959
rect 1719 8956 1731 8959
rect 1762 8956 1768 8968
rect 1719 8928 1768 8956
rect 1719 8925 1731 8928
rect 1673 8919 1731 8925
rect 1762 8916 1768 8928
rect 1820 8956 1826 8968
rect 2317 8959 2375 8965
rect 2317 8956 2329 8959
rect 1820 8928 2329 8956
rect 1820 8916 1826 8928
rect 2317 8925 2329 8928
rect 2363 8925 2375 8959
rect 2317 8919 2375 8925
rect 2406 8916 2412 8968
rect 2464 8916 2470 8968
rect 2608 8965 2636 9120
rect 3142 9092 3148 9104
rect 2700 9064 3148 9092
rect 2700 8965 2728 9064
rect 3142 9052 3148 9064
rect 3200 9092 3206 9104
rect 3970 9092 3976 9104
rect 3200 9064 3976 9092
rect 3200 9052 3206 9064
rect 3970 9052 3976 9064
rect 4028 9052 4034 9104
rect 4080 9092 4108 9132
rect 4341 9129 4353 9163
rect 4387 9160 4399 9163
rect 4706 9160 4712 9172
rect 4387 9132 4712 9160
rect 4387 9129 4399 9132
rect 4341 9123 4399 9129
rect 4706 9120 4712 9132
rect 4764 9120 4770 9172
rect 4890 9120 4896 9172
rect 4948 9160 4954 9172
rect 5534 9160 5540 9172
rect 4948 9132 5540 9160
rect 4948 9120 4954 9132
rect 5534 9120 5540 9132
rect 5592 9120 5598 9172
rect 5810 9120 5816 9172
rect 5868 9120 5874 9172
rect 8570 9120 8576 9172
rect 8628 9120 8634 9172
rect 4080 9064 4568 9092
rect 4540 9024 4568 9064
rect 4982 9052 4988 9104
rect 5040 9092 5046 9104
rect 5040 9064 5856 9092
rect 5040 9052 5046 9064
rect 5828 9024 5856 9064
rect 6914 9052 6920 9104
rect 6972 9092 6978 9104
rect 7834 9092 7840 9104
rect 6972 9064 7840 9092
rect 6972 9052 6978 9064
rect 7834 9052 7840 9064
rect 7892 9052 7898 9104
rect 8297 9095 8355 9101
rect 8297 9061 8309 9095
rect 8343 9092 8355 9095
rect 8588 9092 8616 9120
rect 8343 9064 8616 9092
rect 8343 9061 8355 9064
rect 8297 9055 8355 9061
rect 7742 9024 7748 9036
rect 3804 8996 4476 9024
rect 4540 8996 5764 9024
rect 5828 8996 7748 9024
rect 3804 8965 3832 8996
rect 2593 8959 2651 8965
rect 2593 8925 2605 8959
rect 2639 8925 2651 8959
rect 2593 8919 2651 8925
rect 2685 8959 2743 8965
rect 2685 8925 2697 8959
rect 2731 8925 2743 8959
rect 3789 8959 3847 8965
rect 3789 8956 3801 8959
rect 2685 8919 2743 8925
rect 3712 8928 3801 8956
rect 3712 8900 3740 8928
rect 3789 8925 3801 8928
rect 3835 8925 3847 8959
rect 3789 8919 3847 8925
rect 4154 8916 4160 8968
rect 4212 8916 4218 8968
rect 4448 8965 4476 8996
rect 4249 8959 4307 8965
rect 4249 8925 4261 8959
rect 4295 8925 4307 8959
rect 4249 8919 4307 8925
rect 4433 8959 4491 8965
rect 4433 8925 4445 8959
rect 4479 8925 4491 8959
rect 4433 8919 4491 8925
rect 3694 8848 3700 8900
rect 3752 8848 3758 8900
rect 3878 8848 3884 8900
rect 3936 8888 3942 8900
rect 3973 8891 4031 8897
rect 3973 8888 3985 8891
rect 3936 8860 3985 8888
rect 3936 8848 3942 8860
rect 3973 8857 3985 8860
rect 4019 8888 4031 8891
rect 4264 8888 4292 8919
rect 5258 8916 5264 8968
rect 5316 8956 5322 8968
rect 5442 8956 5448 8968
rect 5316 8928 5448 8956
rect 5316 8916 5322 8928
rect 5442 8916 5448 8928
rect 5500 8956 5506 8968
rect 5736 8966 5764 8996
rect 7742 8984 7748 8996
rect 7800 8984 7806 9036
rect 8018 8984 8024 9036
rect 8076 8984 8082 9036
rect 5537 8959 5595 8965
rect 5537 8956 5549 8959
rect 5500 8928 5549 8956
rect 5500 8916 5506 8928
rect 5537 8925 5549 8928
rect 5583 8925 5595 8959
rect 5736 8938 5856 8966
rect 5537 8919 5595 8925
rect 4019 8860 4292 8888
rect 5552 8888 5580 8919
rect 5828 8897 5856 8938
rect 6914 8916 6920 8968
rect 6972 8916 6978 8968
rect 7926 8916 7932 8968
rect 7984 8916 7990 8968
rect 8757 8959 8815 8965
rect 8757 8925 8769 8959
rect 8803 8956 8815 8959
rect 9306 8956 9312 8968
rect 8803 8928 9312 8956
rect 8803 8925 8815 8928
rect 8757 8919 8815 8925
rect 9306 8916 9312 8928
rect 9364 8916 9370 8968
rect 5813 8891 5871 8897
rect 5552 8860 5764 8888
rect 4019 8857 4031 8860
rect 3973 8851 4031 8857
rect 5166 8780 5172 8832
rect 5224 8820 5230 8832
rect 5629 8823 5687 8829
rect 5629 8820 5641 8823
rect 5224 8792 5641 8820
rect 5224 8780 5230 8792
rect 5629 8789 5641 8792
rect 5675 8789 5687 8823
rect 5736 8820 5764 8860
rect 5813 8857 5825 8891
rect 5859 8888 5871 8891
rect 6932 8888 6960 8916
rect 5859 8860 6960 8888
rect 5859 8857 5871 8860
rect 5813 8851 5871 8857
rect 5994 8820 6000 8832
rect 5736 8792 6000 8820
rect 5629 8783 5687 8789
rect 5994 8780 6000 8792
rect 6052 8820 6058 8832
rect 8573 8823 8631 8829
rect 8573 8820 8585 8823
rect 6052 8792 8585 8820
rect 6052 8780 6058 8792
rect 8573 8789 8585 8792
rect 8619 8789 8631 8823
rect 8573 8783 8631 8789
rect 1104 8730 9384 8752
rect 1104 8678 2645 8730
rect 2697 8678 2709 8730
rect 2761 8678 2773 8730
rect 2825 8678 2837 8730
rect 2889 8678 2901 8730
rect 2953 8678 4715 8730
rect 4767 8678 4779 8730
rect 4831 8678 4843 8730
rect 4895 8678 4907 8730
rect 4959 8678 4971 8730
rect 5023 8678 6785 8730
rect 6837 8678 6849 8730
rect 6901 8678 6913 8730
rect 6965 8678 6977 8730
rect 7029 8678 7041 8730
rect 7093 8678 8855 8730
rect 8907 8678 8919 8730
rect 8971 8678 8983 8730
rect 9035 8678 9047 8730
rect 9099 8678 9111 8730
rect 9163 8678 9384 8730
rect 1104 8656 9384 8678
rect 2225 8619 2283 8625
rect 2225 8585 2237 8619
rect 2271 8616 2283 8619
rect 3694 8616 3700 8628
rect 2271 8588 3700 8616
rect 2271 8585 2283 8588
rect 2225 8579 2283 8585
rect 3694 8576 3700 8588
rect 3752 8616 3758 8628
rect 5166 8616 5172 8628
rect 3752 8588 4200 8616
rect 3752 8576 3758 8588
rect 2406 8548 2412 8560
rect 1872 8520 2412 8548
rect 1872 8489 1900 8520
rect 2406 8508 2412 8520
rect 2464 8548 2470 8560
rect 3050 8548 3056 8560
rect 2464 8520 3056 8548
rect 2464 8508 2470 8520
rect 3050 8508 3056 8520
rect 3108 8508 3114 8560
rect 3878 8508 3884 8560
rect 3936 8548 3942 8560
rect 4172 8557 4200 8588
rect 4264 8588 5172 8616
rect 4264 8557 4292 8588
rect 5166 8576 5172 8588
rect 5224 8576 5230 8628
rect 5261 8619 5319 8625
rect 5261 8585 5273 8619
rect 5307 8616 5319 8619
rect 5350 8616 5356 8628
rect 5307 8588 5356 8616
rect 5307 8585 5319 8588
rect 5261 8579 5319 8585
rect 5350 8576 5356 8588
rect 5408 8576 5414 8628
rect 6914 8576 6920 8628
rect 6972 8616 6978 8628
rect 7101 8619 7159 8625
rect 7101 8616 7113 8619
rect 6972 8588 7113 8616
rect 6972 8576 6978 8588
rect 7101 8585 7113 8588
rect 7147 8616 7159 8619
rect 7558 8616 7564 8628
rect 7147 8588 7564 8616
rect 7147 8585 7159 8588
rect 7101 8579 7159 8585
rect 7558 8576 7564 8588
rect 7616 8576 7622 8628
rect 7926 8576 7932 8628
rect 7984 8616 7990 8628
rect 8297 8619 8355 8625
rect 8297 8616 8309 8619
rect 7984 8588 8309 8616
rect 7984 8576 7990 8588
rect 8297 8585 8309 8588
rect 8343 8585 8355 8619
rect 8297 8579 8355 8585
rect 4157 8551 4215 8557
rect 3936 8520 4016 8548
rect 3936 8508 3942 8520
rect 3988 8489 4016 8520
rect 4157 8517 4169 8551
rect 4203 8517 4215 8551
rect 4157 8511 4215 8517
rect 4249 8551 4307 8557
rect 4249 8517 4261 8551
rect 4295 8517 4307 8551
rect 4249 8511 4307 8517
rect 6733 8551 6791 8557
rect 6733 8517 6745 8551
rect 6779 8548 6791 8551
rect 7653 8551 7711 8557
rect 7653 8548 7665 8551
rect 6779 8520 7665 8548
rect 6779 8517 6791 8520
rect 6733 8511 6791 8517
rect 7653 8517 7665 8520
rect 7699 8548 7711 8551
rect 7699 8520 7880 8548
rect 7699 8517 7711 8520
rect 7653 8511 7711 8517
rect 1857 8483 1915 8489
rect 1857 8449 1869 8483
rect 1903 8449 1915 8483
rect 2961 8483 3019 8489
rect 2961 8480 2973 8483
rect 1857 8443 1915 8449
rect 2424 8452 2973 8480
rect 1762 8372 1768 8424
rect 1820 8372 1826 8424
rect 2424 8288 2452 8452
rect 2961 8449 2973 8452
rect 3007 8449 3019 8483
rect 2961 8443 3019 8449
rect 3973 8483 4031 8489
rect 3973 8449 3985 8483
rect 4019 8449 4031 8483
rect 3973 8443 4031 8449
rect 4341 8483 4399 8489
rect 4341 8449 4353 8483
rect 4387 8480 4399 8483
rect 4430 8480 4436 8492
rect 4387 8452 4436 8480
rect 4387 8449 4399 8452
rect 4341 8443 4399 8449
rect 4430 8440 4436 8452
rect 4488 8440 4494 8492
rect 5169 8483 5227 8489
rect 5169 8449 5181 8483
rect 5215 8480 5227 8483
rect 5258 8480 5264 8492
rect 5215 8452 5264 8480
rect 5215 8449 5227 8452
rect 5169 8443 5227 8449
rect 5258 8440 5264 8452
rect 5316 8440 5322 8492
rect 5350 8440 5356 8492
rect 5408 8440 5414 8492
rect 6917 8483 6975 8489
rect 6917 8449 6929 8483
rect 6963 8480 6975 8483
rect 7006 8480 7012 8492
rect 6963 8452 7012 8480
rect 6963 8449 6975 8452
rect 6917 8443 6975 8449
rect 7006 8440 7012 8452
rect 7064 8440 7070 8492
rect 7190 8440 7196 8492
rect 7248 8440 7254 8492
rect 7852 8489 7880 8520
rect 7469 8483 7527 8489
rect 7469 8449 7481 8483
rect 7515 8480 7527 8483
rect 7745 8483 7803 8489
rect 7515 8452 7604 8480
rect 7515 8449 7527 8452
rect 7469 8443 7527 8449
rect 3237 8415 3295 8421
rect 3237 8381 3249 8415
rect 3283 8412 3295 8415
rect 3510 8412 3516 8424
rect 3283 8384 3516 8412
rect 3283 8381 3295 8384
rect 3237 8375 3295 8381
rect 3510 8372 3516 8384
rect 3568 8372 3574 8424
rect 4522 8304 4528 8356
rect 4580 8304 4586 8356
rect 5994 8304 6000 8356
rect 6052 8344 6058 8356
rect 7285 8347 7343 8353
rect 7285 8344 7297 8347
rect 6052 8316 7297 8344
rect 6052 8304 6058 8316
rect 7285 8313 7297 8316
rect 7331 8313 7343 8347
rect 7285 8307 7343 8313
rect 7576 8288 7604 8452
rect 7745 8449 7757 8483
rect 7791 8449 7803 8483
rect 7745 8443 7803 8449
rect 7837 8483 7895 8489
rect 7837 8449 7849 8483
rect 7883 8449 7895 8483
rect 7837 8443 7895 8449
rect 7760 8412 7788 8443
rect 8662 8440 8668 8492
rect 8720 8440 8726 8492
rect 8018 8412 8024 8424
rect 7760 8384 8024 8412
rect 8018 8372 8024 8384
rect 8076 8372 8082 8424
rect 8941 8347 8999 8353
rect 8941 8313 8953 8347
rect 8987 8344 8999 8347
rect 9030 8344 9036 8356
rect 8987 8316 9036 8344
rect 8987 8313 8999 8316
rect 8941 8307 8999 8313
rect 9030 8304 9036 8316
rect 9088 8304 9094 8356
rect 2406 8236 2412 8288
rect 2464 8236 2470 8288
rect 2774 8236 2780 8288
rect 2832 8236 2838 8288
rect 3145 8279 3203 8285
rect 3145 8245 3157 8279
rect 3191 8276 3203 8279
rect 3234 8276 3240 8288
rect 3191 8248 3240 8276
rect 3191 8245 3203 8248
rect 3145 8239 3203 8245
rect 3234 8236 3240 8248
rect 3292 8276 3298 8288
rect 5902 8276 5908 8288
rect 3292 8248 5908 8276
rect 3292 8236 3298 8248
rect 5902 8236 5908 8248
rect 5960 8236 5966 8288
rect 7558 8236 7564 8288
rect 7616 8276 7622 8288
rect 7929 8279 7987 8285
rect 7929 8276 7941 8279
rect 7616 8248 7941 8276
rect 7616 8236 7622 8248
rect 7929 8245 7941 8248
rect 7975 8245 7987 8279
rect 7929 8239 7987 8245
rect 1104 8186 9384 8208
rect 1104 8134 1985 8186
rect 2037 8134 2049 8186
rect 2101 8134 2113 8186
rect 2165 8134 2177 8186
rect 2229 8134 2241 8186
rect 2293 8134 4055 8186
rect 4107 8134 4119 8186
rect 4171 8134 4183 8186
rect 4235 8134 4247 8186
rect 4299 8134 4311 8186
rect 4363 8134 6125 8186
rect 6177 8134 6189 8186
rect 6241 8134 6253 8186
rect 6305 8134 6317 8186
rect 6369 8134 6381 8186
rect 6433 8134 8195 8186
rect 8247 8134 8259 8186
rect 8311 8134 8323 8186
rect 8375 8134 8387 8186
rect 8439 8134 8451 8186
rect 8503 8134 9384 8186
rect 1104 8112 9384 8134
rect 1762 8032 1768 8084
rect 1820 8072 1826 8084
rect 1949 8075 2007 8081
rect 1949 8072 1961 8075
rect 1820 8044 1961 8072
rect 1820 8032 1826 8044
rect 1949 8041 1961 8044
rect 1995 8041 2007 8075
rect 1949 8035 2007 8041
rect 5074 8032 5080 8084
rect 5132 8032 5138 8084
rect 5442 8072 5448 8084
rect 5184 8044 5448 8072
rect 5184 8004 5212 8044
rect 5442 8032 5448 8044
rect 5500 8032 5506 8084
rect 6914 8032 6920 8084
rect 6972 8032 6978 8084
rect 7190 8032 7196 8084
rect 7248 8072 7254 8084
rect 7374 8072 7380 8084
rect 7248 8044 7380 8072
rect 7248 8032 7254 8044
rect 7374 8032 7380 8044
rect 7432 8072 7438 8084
rect 7469 8075 7527 8081
rect 7469 8072 7481 8075
rect 7432 8044 7481 8072
rect 7432 8032 7438 8044
rect 7469 8041 7481 8044
rect 7515 8041 7527 8075
rect 7469 8035 7527 8041
rect 7558 8032 7564 8084
rect 7616 8032 7622 8084
rect 7650 8032 7656 8084
rect 7708 8072 7714 8084
rect 7745 8075 7803 8081
rect 7745 8072 7757 8075
rect 7708 8044 7757 8072
rect 7708 8032 7714 8044
rect 7745 8041 7757 8044
rect 7791 8041 7803 8075
rect 7745 8035 7803 8041
rect 8018 8032 8024 8084
rect 8076 8032 8082 8084
rect 8389 8075 8447 8081
rect 8389 8041 8401 8075
rect 8435 8072 8447 8075
rect 8570 8072 8576 8084
rect 8435 8044 8576 8072
rect 8435 8041 8447 8044
rect 8389 8035 8447 8041
rect 8570 8032 8576 8044
rect 8628 8032 8634 8084
rect 3528 7976 5212 8004
rect 2685 7939 2743 7945
rect 2685 7936 2697 7939
rect 2148 7908 2697 7936
rect 2148 7877 2176 7908
rect 2685 7905 2697 7908
rect 2731 7936 2743 7939
rect 2774 7936 2780 7948
rect 2731 7908 2780 7936
rect 2731 7905 2743 7908
rect 2685 7899 2743 7905
rect 2774 7896 2780 7908
rect 2832 7896 2838 7948
rect 2133 7871 2191 7877
rect 2133 7837 2145 7871
rect 2179 7837 2191 7871
rect 2133 7831 2191 7837
rect 2406 7828 2412 7880
rect 2464 7828 2470 7880
rect 2961 7871 3019 7877
rect 2961 7868 2973 7871
rect 2700 7840 2973 7868
rect 2314 7760 2320 7812
rect 2372 7800 2378 7812
rect 2700 7800 2728 7840
rect 2961 7837 2973 7840
rect 3007 7868 3019 7871
rect 3528 7868 3556 7976
rect 5258 7964 5264 8016
rect 5316 8004 5322 8016
rect 5629 8007 5687 8013
rect 5629 8004 5641 8007
rect 5316 7976 5641 8004
rect 5316 7964 5322 7976
rect 5629 7973 5641 7976
rect 5675 7973 5687 8007
rect 5629 7967 5687 7973
rect 3605 7939 3663 7945
rect 3605 7905 3617 7939
rect 3651 7936 3663 7939
rect 4430 7936 4436 7948
rect 3651 7908 4436 7936
rect 3651 7905 3663 7908
rect 3605 7899 3663 7905
rect 4430 7896 4436 7908
rect 4488 7936 4494 7948
rect 4525 7939 4583 7945
rect 4525 7936 4537 7939
rect 4488 7908 4537 7936
rect 4488 7896 4494 7908
rect 4525 7905 4537 7908
rect 4571 7905 4583 7939
rect 4525 7899 4583 7905
rect 4985 7939 5043 7945
rect 4985 7905 4997 7939
rect 5031 7936 5043 7939
rect 5442 7936 5448 7948
rect 5031 7908 5448 7936
rect 5031 7905 5043 7908
rect 4985 7899 5043 7905
rect 3007 7840 3556 7868
rect 3007 7837 3019 7840
rect 2961 7831 3019 7837
rect 2372 7772 2728 7800
rect 4540 7800 4568 7899
rect 5442 7896 5448 7908
rect 5500 7936 5506 7948
rect 5500 7908 5856 7936
rect 5500 7896 5506 7908
rect 4617 7871 4675 7877
rect 4617 7837 4629 7871
rect 4663 7868 4675 7871
rect 5166 7868 5172 7880
rect 4663 7840 5172 7868
rect 4663 7837 4675 7840
rect 4617 7831 4675 7837
rect 5166 7828 5172 7840
rect 5224 7828 5230 7880
rect 5258 7828 5264 7880
rect 5316 7828 5322 7880
rect 5828 7877 5856 7908
rect 5902 7896 5908 7948
rect 5960 7896 5966 7948
rect 5994 7896 6000 7948
rect 6052 7896 6058 7948
rect 6288 7908 6868 7936
rect 5537 7871 5595 7877
rect 5537 7837 5549 7871
rect 5583 7837 5595 7871
rect 5537 7831 5595 7837
rect 5813 7871 5871 7877
rect 5813 7837 5825 7871
rect 5859 7837 5871 7871
rect 5920 7868 5948 7896
rect 6288 7877 6316 7908
rect 6273 7871 6331 7877
rect 6273 7868 6285 7871
rect 5920 7840 6285 7868
rect 5813 7831 5871 7837
rect 6273 7837 6285 7840
rect 6319 7837 6331 7871
rect 6273 7831 6331 7837
rect 5552 7800 5580 7831
rect 6362 7828 6368 7880
rect 6420 7868 6426 7880
rect 6641 7871 6699 7877
rect 6641 7868 6653 7871
rect 6420 7840 6653 7868
rect 6420 7828 6426 7840
rect 6641 7837 6653 7840
rect 6687 7837 6699 7871
rect 6641 7831 6699 7837
rect 6733 7871 6791 7877
rect 6733 7837 6745 7871
rect 6779 7837 6791 7871
rect 6840 7868 6868 7908
rect 7083 7871 7141 7877
rect 6840 7862 6960 7868
rect 7083 7862 7095 7871
rect 6840 7840 7095 7862
rect 6733 7831 6791 7837
rect 6932 7837 7095 7840
rect 7129 7837 7141 7871
rect 6932 7834 7141 7837
rect 7083 7831 7141 7834
rect 4540 7772 5580 7800
rect 2372 7760 2378 7772
rect 6086 7760 6092 7812
rect 6144 7800 6150 7812
rect 6757 7800 6785 7831
rect 7190 7828 7196 7880
rect 7248 7828 7254 7880
rect 7285 7871 7343 7877
rect 7285 7837 7297 7871
rect 7331 7837 7343 7871
rect 7285 7831 7343 7837
rect 7300 7800 7328 7831
rect 7374 7828 7380 7880
rect 7432 7828 7438 7880
rect 8481 7871 8539 7877
rect 8481 7837 8493 7871
rect 8527 7837 8539 7871
rect 8481 7831 8539 7837
rect 6144 7772 7328 7800
rect 7392 7800 7420 7828
rect 7713 7803 7771 7809
rect 7713 7800 7725 7803
rect 7392 7772 7725 7800
rect 6144 7760 6150 7772
rect 7713 7769 7725 7772
rect 7759 7769 7771 7803
rect 7713 7763 7771 7769
rect 7929 7803 7987 7809
rect 7929 7769 7941 7803
rect 7975 7800 7987 7803
rect 8110 7800 8116 7812
rect 7975 7772 8116 7800
rect 7975 7769 7987 7772
rect 7929 7763 7987 7769
rect 5166 7692 5172 7744
rect 5224 7732 5230 7744
rect 5445 7735 5503 7741
rect 5445 7732 5457 7735
rect 5224 7704 5457 7732
rect 5224 7692 5230 7704
rect 5445 7701 5457 7704
rect 5491 7732 5503 7735
rect 5902 7732 5908 7744
rect 5491 7704 5908 7732
rect 5491 7701 5503 7704
rect 5445 7695 5503 7701
rect 5902 7692 5908 7704
rect 5960 7692 5966 7744
rect 7006 7692 7012 7744
rect 7064 7732 7070 7744
rect 7944 7732 7972 7763
rect 8110 7760 8116 7772
rect 8168 7760 8174 7812
rect 8496 7744 8524 7831
rect 7064 7704 7972 7732
rect 7064 7692 7070 7704
rect 8478 7692 8484 7744
rect 8536 7692 8542 7744
rect 1104 7642 9384 7664
rect 1104 7590 2645 7642
rect 2697 7590 2709 7642
rect 2761 7590 2773 7642
rect 2825 7590 2837 7642
rect 2889 7590 2901 7642
rect 2953 7590 4715 7642
rect 4767 7590 4779 7642
rect 4831 7590 4843 7642
rect 4895 7590 4907 7642
rect 4959 7590 4971 7642
rect 5023 7590 6785 7642
rect 6837 7590 6849 7642
rect 6901 7590 6913 7642
rect 6965 7590 6977 7642
rect 7029 7590 7041 7642
rect 7093 7590 8855 7642
rect 8907 7590 8919 7642
rect 8971 7590 8983 7642
rect 9035 7590 9047 7642
rect 9099 7590 9111 7642
rect 9163 7590 9384 7642
rect 1104 7568 9384 7590
rect 2314 7488 2320 7540
rect 2372 7528 2378 7540
rect 5261 7531 5319 7537
rect 2372 7500 2774 7528
rect 2372 7488 2378 7500
rect 2746 7460 2774 7500
rect 5261 7497 5273 7531
rect 5307 7528 5319 7531
rect 5350 7528 5356 7540
rect 5307 7500 5356 7528
rect 5307 7497 5319 7500
rect 5261 7491 5319 7497
rect 5350 7488 5356 7500
rect 5408 7488 5414 7540
rect 5442 7488 5448 7540
rect 5500 7488 5506 7540
rect 5994 7488 6000 7540
rect 6052 7488 6058 7540
rect 8662 7488 8668 7540
rect 8720 7528 8726 7540
rect 8849 7531 8907 7537
rect 8849 7528 8861 7531
rect 8720 7500 8861 7528
rect 8720 7488 8726 7500
rect 8849 7497 8861 7500
rect 8895 7497 8907 7531
rect 8849 7491 8907 7497
rect 2746 7432 2912 7460
rect 1762 7352 1768 7404
rect 1820 7352 1826 7404
rect 2406 7352 2412 7404
rect 2464 7392 2470 7404
rect 2682 7392 2688 7404
rect 2464 7364 2688 7392
rect 2464 7352 2470 7364
rect 2682 7352 2688 7364
rect 2740 7352 2746 7404
rect 2884 7401 2912 7432
rect 2869 7395 2927 7401
rect 2869 7361 2881 7395
rect 2915 7361 2927 7395
rect 2869 7355 2927 7361
rect 3145 7395 3203 7401
rect 3145 7361 3157 7395
rect 3191 7392 3203 7395
rect 3510 7392 3516 7404
rect 3191 7364 3516 7392
rect 3191 7361 3203 7364
rect 3145 7355 3203 7361
rect 3510 7352 3516 7364
rect 3568 7392 3574 7404
rect 5460 7401 5488 7488
rect 5445 7395 5503 7401
rect 3568 7364 5396 7392
rect 3568 7352 3574 7364
rect 2961 7327 3019 7333
rect 2961 7293 2973 7327
rect 3007 7324 3019 7327
rect 3234 7324 3240 7336
rect 3007 7296 3240 7324
rect 3007 7293 3019 7296
rect 2961 7287 3019 7293
rect 3234 7284 3240 7296
rect 3292 7284 3298 7336
rect 5261 7327 5319 7333
rect 5261 7324 5273 7327
rect 5184 7296 5273 7324
rect 2777 7259 2835 7265
rect 2777 7225 2789 7259
rect 2823 7256 2835 7259
rect 5184 7256 5212 7296
rect 5261 7293 5273 7296
rect 5307 7293 5319 7327
rect 5368 7324 5396 7364
rect 5445 7361 5457 7395
rect 5491 7361 5503 7395
rect 5445 7355 5503 7361
rect 5537 7395 5595 7401
rect 5537 7361 5549 7395
rect 5583 7392 5595 7395
rect 6012 7392 6040 7488
rect 5583 7364 6040 7392
rect 5583 7361 5595 7364
rect 5537 7355 5595 7361
rect 8662 7352 8668 7404
rect 8720 7352 8726 7404
rect 6362 7324 6368 7336
rect 5368 7296 6368 7324
rect 5261 7287 5319 7293
rect 6362 7284 6368 7296
rect 6420 7324 6426 7336
rect 7190 7324 7196 7336
rect 6420 7296 7196 7324
rect 6420 7284 6426 7296
rect 7190 7284 7196 7296
rect 7248 7284 7254 7336
rect 8389 7327 8447 7333
rect 8389 7293 8401 7327
rect 8435 7324 8447 7327
rect 8570 7324 8576 7336
rect 8435 7296 8576 7324
rect 8435 7293 8447 7296
rect 8389 7287 8447 7293
rect 8570 7284 8576 7296
rect 8628 7284 8634 7336
rect 5534 7256 5540 7268
rect 2823 7228 3096 7256
rect 2823 7225 2835 7228
rect 2777 7219 2835 7225
rect 3068 7200 3096 7228
rect 5184 7228 5540 7256
rect 5184 7200 5212 7228
rect 5534 7216 5540 7228
rect 5592 7216 5598 7268
rect 7208 7256 7236 7284
rect 8018 7256 8024 7268
rect 7208 7228 8024 7256
rect 8018 7216 8024 7228
rect 8076 7256 8082 7268
rect 8478 7256 8484 7268
rect 8076 7228 8484 7256
rect 8076 7216 8082 7228
rect 8478 7216 8484 7228
rect 8536 7216 8542 7268
rect 1486 7148 1492 7200
rect 1544 7148 1550 7200
rect 2406 7148 2412 7200
rect 2464 7148 2470 7200
rect 3050 7148 3056 7200
rect 3108 7148 3114 7200
rect 5166 7148 5172 7200
rect 5224 7148 5230 7200
rect 1104 7098 9384 7120
rect 1104 7046 1985 7098
rect 2037 7046 2049 7098
rect 2101 7046 2113 7098
rect 2165 7046 2177 7098
rect 2229 7046 2241 7098
rect 2293 7046 4055 7098
rect 4107 7046 4119 7098
rect 4171 7046 4183 7098
rect 4235 7046 4247 7098
rect 4299 7046 4311 7098
rect 4363 7046 6125 7098
rect 6177 7046 6189 7098
rect 6241 7046 6253 7098
rect 6305 7046 6317 7098
rect 6369 7046 6381 7098
rect 6433 7046 8195 7098
rect 8247 7046 8259 7098
rect 8311 7046 8323 7098
rect 8375 7046 8387 7098
rect 8439 7046 8451 7098
rect 8503 7046 9384 7098
rect 1104 7024 9384 7046
rect 2130 6944 2136 6996
rect 2188 6984 2194 6996
rect 2682 6984 2688 6996
rect 2188 6956 2688 6984
rect 2188 6944 2194 6956
rect 2682 6944 2688 6956
rect 2740 6984 2746 6996
rect 4706 6984 4712 6996
rect 2740 6956 4712 6984
rect 2740 6944 2746 6956
rect 4706 6944 4712 6956
rect 4764 6984 4770 6996
rect 5994 6984 6000 6996
rect 4764 6956 6000 6984
rect 4764 6944 4770 6956
rect 5994 6944 6000 6956
rect 6052 6944 6058 6996
rect 1780 6888 2452 6916
rect 1780 6857 1808 6888
rect 2424 6860 2452 6888
rect 7374 6876 7380 6928
rect 7432 6916 7438 6928
rect 7742 6916 7748 6928
rect 7432 6888 7748 6916
rect 7432 6876 7438 6888
rect 7742 6876 7748 6888
rect 7800 6916 7806 6928
rect 7929 6919 7987 6925
rect 7929 6916 7941 6919
rect 7800 6888 7941 6916
rect 7800 6876 7806 6888
rect 7929 6885 7941 6888
rect 7975 6885 7987 6919
rect 7929 6879 7987 6885
rect 8018 6876 8024 6928
rect 8076 6876 8082 6928
rect 1765 6851 1823 6857
rect 1765 6817 1777 6851
rect 1811 6848 1823 6851
rect 2041 6851 2099 6857
rect 1811 6820 1845 6848
rect 1811 6817 1823 6820
rect 1765 6811 1823 6817
rect 2041 6817 2053 6851
rect 2087 6848 2099 6851
rect 2314 6848 2320 6860
rect 2087 6820 2320 6848
rect 2087 6817 2099 6820
rect 2041 6811 2099 6817
rect 2314 6808 2320 6820
rect 2372 6808 2378 6860
rect 2406 6808 2412 6860
rect 2464 6808 2470 6860
rect 3789 6851 3847 6857
rect 3789 6817 3801 6851
rect 3835 6848 3847 6851
rect 4154 6848 4160 6860
rect 3835 6820 4160 6848
rect 3835 6817 3847 6820
rect 3789 6811 3847 6817
rect 4154 6808 4160 6820
rect 4212 6848 4218 6860
rect 4614 6848 4620 6860
rect 4212 6820 4620 6848
rect 4212 6808 4218 6820
rect 4614 6808 4620 6820
rect 4672 6808 4678 6860
rect 6656 6820 7696 6848
rect 6656 6792 6684 6820
rect 7668 6792 7696 6820
rect 1673 6783 1731 6789
rect 1673 6749 1685 6783
rect 1719 6780 1731 6783
rect 1854 6780 1860 6792
rect 1719 6752 1860 6780
rect 1719 6749 1731 6752
rect 1673 6743 1731 6749
rect 1854 6740 1860 6752
rect 1912 6740 1918 6792
rect 3973 6783 4031 6789
rect 3973 6749 3985 6783
rect 4019 6749 4031 6783
rect 3973 6743 4031 6749
rect 4341 6783 4399 6789
rect 4341 6749 4353 6783
rect 4387 6780 4399 6783
rect 4522 6780 4528 6792
rect 4387 6752 4528 6780
rect 4387 6749 4399 6752
rect 4341 6743 4399 6749
rect 3878 6672 3884 6724
rect 3936 6672 3942 6724
rect 3988 6656 4016 6743
rect 4522 6740 4528 6752
rect 4580 6740 4586 6792
rect 6638 6740 6644 6792
rect 6696 6740 6702 6792
rect 7190 6740 7196 6792
rect 7248 6780 7254 6792
rect 7285 6783 7343 6789
rect 7285 6780 7297 6783
rect 7248 6752 7297 6780
rect 7248 6740 7254 6752
rect 7285 6749 7297 6752
rect 7331 6749 7343 6783
rect 7285 6743 7343 6749
rect 7650 6740 7656 6792
rect 7708 6740 7714 6792
rect 7926 6740 7932 6792
rect 7984 6740 7990 6792
rect 8036 6780 8064 6876
rect 8386 6780 8392 6792
rect 8036 6752 8392 6780
rect 8386 6740 8392 6752
rect 8444 6740 8450 6792
rect 4617 6715 4675 6721
rect 4617 6681 4629 6715
rect 4663 6712 4675 6715
rect 5258 6712 5264 6724
rect 4663 6684 5264 6712
rect 4663 6681 4675 6684
rect 4617 6675 4675 6681
rect 3970 6604 3976 6656
rect 4028 6604 4034 6656
rect 4338 6604 4344 6656
rect 4396 6644 4402 6656
rect 4632 6644 4660 6675
rect 5258 6672 5264 6684
rect 5316 6672 5322 6724
rect 7668 6712 7696 6740
rect 8113 6715 8171 6721
rect 8113 6712 8125 6715
rect 7668 6684 8125 6712
rect 8113 6681 8125 6684
rect 8159 6681 8171 6715
rect 8113 6675 8171 6681
rect 4396 6616 4660 6644
rect 7469 6647 7527 6653
rect 4396 6604 4402 6616
rect 7469 6613 7481 6647
rect 7515 6644 7527 6647
rect 7834 6644 7840 6656
rect 7515 6616 7840 6644
rect 7515 6613 7527 6616
rect 7469 6607 7527 6613
rect 7834 6604 7840 6616
rect 7892 6604 7898 6656
rect 8202 6604 8208 6656
rect 8260 6653 8266 6656
rect 8260 6607 8269 6653
rect 8297 6647 8355 6653
rect 8297 6613 8309 6647
rect 8343 6644 8355 6647
rect 8478 6644 8484 6656
rect 8343 6616 8484 6644
rect 8343 6613 8355 6616
rect 8297 6607 8355 6613
rect 8260 6604 8266 6607
rect 8478 6604 8484 6616
rect 8536 6604 8542 6656
rect 1104 6554 9384 6576
rect 1104 6502 2645 6554
rect 2697 6502 2709 6554
rect 2761 6502 2773 6554
rect 2825 6502 2837 6554
rect 2889 6502 2901 6554
rect 2953 6502 4715 6554
rect 4767 6502 4779 6554
rect 4831 6502 4843 6554
rect 4895 6502 4907 6554
rect 4959 6502 4971 6554
rect 5023 6502 6785 6554
rect 6837 6502 6849 6554
rect 6901 6502 6913 6554
rect 6965 6502 6977 6554
rect 7029 6502 7041 6554
rect 7093 6502 8855 6554
rect 8907 6502 8919 6554
rect 8971 6502 8983 6554
rect 9035 6502 9047 6554
rect 9099 6502 9111 6554
rect 9163 6502 9384 6554
rect 1104 6480 9384 6502
rect 1854 6400 1860 6452
rect 1912 6440 1918 6452
rect 2225 6443 2283 6449
rect 2225 6440 2237 6443
rect 1912 6412 2237 6440
rect 1912 6400 1918 6412
rect 2225 6409 2237 6412
rect 2271 6409 2283 6443
rect 2225 6403 2283 6409
rect 4338 6400 4344 6452
rect 4396 6440 4402 6452
rect 4396 6412 4844 6440
rect 4396 6400 4402 6412
rect 2130 6332 2136 6384
rect 2188 6332 2194 6384
rect 2593 6375 2651 6381
rect 2593 6341 2605 6375
rect 2639 6372 2651 6375
rect 3234 6372 3240 6384
rect 2639 6344 3240 6372
rect 2639 6341 2651 6344
rect 2593 6335 2651 6341
rect 3234 6332 3240 6344
rect 3292 6332 3298 6384
rect 3970 6372 3976 6384
rect 3620 6344 3976 6372
rect 2136 6329 2194 6332
rect 2136 6295 2148 6329
rect 2182 6295 2194 6329
rect 2136 6289 2194 6295
rect 2406 6264 2412 6316
rect 2464 6264 2470 6316
rect 3620 6313 3648 6344
rect 3970 6332 3976 6344
rect 4028 6372 4034 6384
rect 4028 6344 4660 6372
rect 4028 6332 4034 6344
rect 3605 6307 3663 6313
rect 3605 6304 3617 6307
rect 2792 6276 3617 6304
rect 2792 6112 2820 6276
rect 3605 6273 3617 6276
rect 3651 6273 3663 6307
rect 3605 6267 3663 6273
rect 3789 6307 3847 6313
rect 3789 6273 3801 6307
rect 3835 6304 3847 6307
rect 3881 6307 3939 6313
rect 3881 6304 3893 6307
rect 3835 6276 3893 6304
rect 3835 6273 3847 6276
rect 3789 6267 3847 6273
rect 3881 6273 3893 6276
rect 3927 6273 3939 6307
rect 3881 6267 3939 6273
rect 4065 6307 4123 6313
rect 4065 6273 4077 6307
rect 4111 6304 4123 6307
rect 4154 6304 4160 6316
rect 4111 6276 4160 6304
rect 4111 6273 4123 6276
rect 4065 6267 4123 6273
rect 4154 6264 4160 6276
rect 4212 6304 4218 6316
rect 4632 6313 4660 6344
rect 4816 6313 4844 6412
rect 5994 6400 6000 6452
rect 6052 6400 6058 6452
rect 7101 6443 7159 6449
rect 7101 6440 7113 6443
rect 6196 6412 7113 6440
rect 6196 6313 6224 6412
rect 7101 6409 7113 6412
rect 7147 6409 7159 6443
rect 7101 6403 7159 6409
rect 7650 6400 7656 6452
rect 7708 6440 7714 6452
rect 7708 6412 8065 6440
rect 7708 6400 7714 6412
rect 6638 6332 6644 6384
rect 6696 6372 6702 6384
rect 6742 6375 6800 6381
rect 6742 6372 6754 6375
rect 6696 6344 6754 6372
rect 6696 6332 6702 6344
rect 6742 6341 6754 6344
rect 6788 6341 6800 6375
rect 6742 6335 6800 6341
rect 7576 6344 7972 6372
rect 7576 6316 7604 6344
rect 4433 6307 4491 6313
rect 4433 6304 4445 6307
rect 4212 6276 4445 6304
rect 4212 6264 4218 6276
rect 4433 6273 4445 6276
rect 4479 6273 4491 6307
rect 4433 6267 4491 6273
rect 4617 6307 4675 6313
rect 4617 6273 4629 6307
rect 4663 6273 4675 6307
rect 4617 6267 4675 6273
rect 4709 6307 4767 6313
rect 4709 6273 4721 6307
rect 4755 6273 4767 6307
rect 4709 6267 4767 6273
rect 4801 6307 4859 6313
rect 4801 6273 4813 6307
rect 4847 6273 4859 6307
rect 4801 6267 4859 6273
rect 6181 6307 6239 6313
rect 6181 6273 6193 6307
rect 6227 6273 6239 6307
rect 6181 6267 6239 6273
rect 6365 6307 6423 6313
rect 6365 6273 6377 6307
rect 6411 6304 6423 6307
rect 7377 6307 7435 6313
rect 7377 6304 7389 6307
rect 6411 6276 7389 6304
rect 6411 6273 6423 6276
rect 6365 6267 6423 6273
rect 7377 6273 7389 6276
rect 7423 6273 7435 6307
rect 7377 6267 7435 6273
rect 4338 6196 4344 6248
rect 4396 6196 4402 6248
rect 4724 6236 4752 6267
rect 4540 6208 4752 6236
rect 7392 6236 7420 6267
rect 7558 6264 7564 6316
rect 7616 6264 7622 6316
rect 7650 6264 7656 6316
rect 7708 6264 7714 6316
rect 7944 6313 7972 6344
rect 8037 6313 8065 6412
rect 8202 6400 8208 6452
rect 8260 6400 8266 6452
rect 8662 6400 8668 6452
rect 8720 6400 8726 6452
rect 8220 6372 8248 6400
rect 8220 6344 8984 6372
rect 7929 6307 7987 6313
rect 7929 6273 7941 6307
rect 7975 6273 7987 6307
rect 7929 6267 7987 6273
rect 8022 6307 8080 6313
rect 8022 6273 8034 6307
rect 8068 6273 8080 6307
rect 8022 6267 8080 6273
rect 8205 6307 8263 6313
rect 8205 6273 8217 6307
rect 8251 6273 8263 6307
rect 8205 6267 8263 6273
rect 8297 6307 8355 6313
rect 8297 6273 8309 6307
rect 8343 6273 8355 6307
rect 8297 6267 8355 6273
rect 8220 6236 8248 6267
rect 7392 6208 8248 6236
rect 8312 6236 8340 6267
rect 8386 6264 8392 6316
rect 8444 6313 8450 6316
rect 8956 6313 8984 6344
rect 8444 6304 8452 6313
rect 8941 6307 8999 6313
rect 8444 6276 8489 6304
rect 8444 6267 8452 6276
rect 8941 6273 8953 6307
rect 8987 6273 8999 6307
rect 8941 6267 8999 6273
rect 8444 6264 8450 6267
rect 8665 6239 8723 6245
rect 8665 6236 8677 6239
rect 8312 6208 8524 6236
rect 4540 6112 4568 6208
rect 6748 6140 7604 6168
rect 2774 6060 2780 6112
rect 2832 6060 2838 6112
rect 3418 6060 3424 6112
rect 3476 6060 3482 6112
rect 4249 6103 4307 6109
rect 4249 6069 4261 6103
rect 4295 6100 4307 6103
rect 4522 6100 4528 6112
rect 4295 6072 4528 6100
rect 4295 6069 4307 6072
rect 4249 6063 4307 6069
rect 4522 6060 4528 6072
rect 4580 6060 4586 6112
rect 5074 6060 5080 6112
rect 5132 6060 5138 6112
rect 6748 6109 6776 6140
rect 7576 6112 7604 6140
rect 7668 6112 7696 6208
rect 8496 6180 8524 6208
rect 8588 6208 8677 6236
rect 7926 6128 7932 6180
rect 7984 6128 7990 6180
rect 8478 6128 8484 6180
rect 8536 6128 8542 6180
rect 8588 6177 8616 6208
rect 8665 6205 8677 6208
rect 8711 6205 8723 6239
rect 8665 6199 8723 6205
rect 8573 6171 8631 6177
rect 8573 6137 8585 6171
rect 8619 6137 8631 6171
rect 8573 6131 8631 6137
rect 6733 6103 6791 6109
rect 6733 6069 6745 6103
rect 6779 6069 6791 6103
rect 6733 6063 6791 6069
rect 6822 6060 6828 6112
rect 6880 6100 6886 6112
rect 6917 6103 6975 6109
rect 6917 6100 6929 6103
rect 6880 6072 6929 6100
rect 6880 6060 6886 6072
rect 6917 6069 6929 6072
rect 6963 6100 6975 6103
rect 7466 6100 7472 6112
rect 6963 6072 7472 6100
rect 6963 6069 6975 6072
rect 6917 6063 6975 6069
rect 7466 6060 7472 6072
rect 7524 6060 7530 6112
rect 7558 6060 7564 6112
rect 7616 6060 7622 6112
rect 7650 6060 7656 6112
rect 7708 6060 7714 6112
rect 7944 6100 7972 6128
rect 8849 6103 8907 6109
rect 8849 6100 8861 6103
rect 7944 6072 8861 6100
rect 8849 6069 8861 6072
rect 8895 6069 8907 6103
rect 8849 6063 8907 6069
rect 1104 6010 9384 6032
rect 1104 5958 1985 6010
rect 2037 5958 2049 6010
rect 2101 5958 2113 6010
rect 2165 5958 2177 6010
rect 2229 5958 2241 6010
rect 2293 5958 4055 6010
rect 4107 5958 4119 6010
rect 4171 5958 4183 6010
rect 4235 5958 4247 6010
rect 4299 5958 4311 6010
rect 4363 5958 6125 6010
rect 6177 5958 6189 6010
rect 6241 5958 6253 6010
rect 6305 5958 6317 6010
rect 6369 5958 6381 6010
rect 6433 5958 8195 6010
rect 8247 5958 8259 6010
rect 8311 5958 8323 6010
rect 8375 5958 8387 6010
rect 8439 5958 8451 6010
rect 8503 5958 9384 6010
rect 1104 5936 9384 5958
rect 1854 5856 1860 5908
rect 1912 5856 1918 5908
rect 2774 5856 2780 5908
rect 2832 5856 2838 5908
rect 3418 5856 3424 5908
rect 3476 5856 3482 5908
rect 4985 5899 5043 5905
rect 4985 5865 4997 5899
rect 5031 5896 5043 5899
rect 5350 5896 5356 5908
rect 5031 5868 5356 5896
rect 5031 5865 5043 5868
rect 4985 5859 5043 5865
rect 5350 5856 5356 5868
rect 5408 5856 5414 5908
rect 6638 5856 6644 5908
rect 6696 5856 6702 5908
rect 7101 5899 7159 5905
rect 7101 5865 7113 5899
rect 7147 5896 7159 5899
rect 7190 5896 7196 5908
rect 7147 5868 7196 5896
rect 7147 5865 7159 5868
rect 7101 5859 7159 5865
rect 7190 5856 7196 5868
rect 7248 5856 7254 5908
rect 7285 5899 7343 5905
rect 7285 5865 7297 5899
rect 7331 5865 7343 5899
rect 7837 5899 7895 5905
rect 7837 5896 7849 5899
rect 7285 5859 7343 5865
rect 7668 5868 7849 5896
rect 1872 5760 1900 5856
rect 2225 5831 2283 5837
rect 2225 5797 2237 5831
rect 2271 5828 2283 5831
rect 3436 5828 3464 5856
rect 6656 5828 6684 5856
rect 7300 5828 7328 5859
rect 2271 5800 2774 5828
rect 3436 5800 4108 5828
rect 6656 5800 7328 5828
rect 2271 5797 2283 5800
rect 2225 5791 2283 5797
rect 1949 5763 2007 5769
rect 1949 5760 1961 5763
rect 1872 5732 1961 5760
rect 1949 5729 1961 5732
rect 1995 5760 2007 5763
rect 2130 5760 2136 5772
rect 1995 5732 2136 5760
rect 1995 5729 2007 5732
rect 1949 5723 2007 5729
rect 2130 5720 2136 5732
rect 2188 5720 2194 5772
rect 2314 5720 2320 5772
rect 2372 5760 2378 5772
rect 2409 5763 2467 5769
rect 2409 5760 2421 5763
rect 2372 5732 2421 5760
rect 2372 5720 2378 5732
rect 2409 5729 2421 5732
rect 2455 5729 2467 5763
rect 2746 5760 2774 5800
rect 3973 5763 4031 5769
rect 3973 5760 3985 5763
rect 2746 5732 3985 5760
rect 2409 5723 2467 5729
rect 3973 5729 3985 5732
rect 4019 5729 4031 5763
rect 4080 5760 4108 5800
rect 4249 5763 4307 5769
rect 4249 5760 4261 5763
rect 4080 5732 4261 5760
rect 3973 5723 4031 5729
rect 4249 5729 4261 5732
rect 4295 5729 4307 5763
rect 4801 5763 4859 5769
rect 4801 5760 4813 5763
rect 4249 5723 4307 5729
rect 4448 5732 4813 5760
rect 4448 5704 4476 5732
rect 4801 5729 4813 5732
rect 4847 5729 4859 5763
rect 4801 5723 4859 5729
rect 7668 5704 7696 5868
rect 7837 5865 7849 5868
rect 7883 5865 7895 5899
rect 7837 5859 7895 5865
rect 7926 5856 7932 5908
rect 7984 5896 7990 5908
rect 8205 5899 8263 5905
rect 8205 5896 8217 5899
rect 7984 5868 8217 5896
rect 7984 5856 7990 5868
rect 8205 5865 8217 5868
rect 8251 5865 8263 5899
rect 8205 5859 8263 5865
rect 8662 5856 8668 5908
rect 8720 5856 8726 5908
rect 1578 5652 1584 5704
rect 1636 5652 1642 5704
rect 1762 5652 1768 5704
rect 1820 5652 1826 5704
rect 1857 5695 1915 5701
rect 1857 5661 1869 5695
rect 1903 5661 1915 5695
rect 1857 5655 1915 5661
rect 2041 5695 2099 5701
rect 2041 5661 2053 5695
rect 2087 5692 2099 5695
rect 2222 5692 2228 5704
rect 2087 5664 2228 5692
rect 2087 5661 2099 5664
rect 2041 5655 2099 5661
rect 1596 5624 1624 5652
rect 1872 5624 1900 5655
rect 2222 5652 2228 5664
rect 2280 5652 2286 5704
rect 2501 5695 2559 5701
rect 2501 5661 2513 5695
rect 2547 5661 2559 5695
rect 2501 5655 2559 5661
rect 2516 5624 2544 5655
rect 3142 5652 3148 5704
rect 3200 5652 3206 5704
rect 3878 5652 3884 5704
rect 3936 5652 3942 5704
rect 4062 5652 4068 5704
rect 4120 5652 4126 5704
rect 4157 5695 4215 5701
rect 4157 5661 4169 5695
rect 4203 5661 4215 5695
rect 4157 5655 4215 5661
rect 1596 5596 2544 5624
rect 1946 5516 1952 5568
rect 2004 5556 2010 5568
rect 3160 5556 3188 5652
rect 3896 5624 3924 5652
rect 4172 5624 4200 5655
rect 4430 5652 4436 5704
rect 4488 5652 4494 5704
rect 5074 5652 5080 5704
rect 5132 5652 5138 5704
rect 7377 5695 7435 5701
rect 7377 5661 7389 5695
rect 7423 5661 7435 5695
rect 7377 5655 7435 5661
rect 5810 5624 5816 5636
rect 3896 5596 4200 5624
rect 4448 5596 5816 5624
rect 4448 5565 4476 5596
rect 5810 5584 5816 5596
rect 5868 5584 5874 5636
rect 7392 5624 7420 5655
rect 7650 5652 7656 5704
rect 7708 5652 7714 5704
rect 7745 5695 7803 5701
rect 7745 5661 7757 5695
rect 7791 5661 7803 5695
rect 7745 5655 7803 5661
rect 7558 5624 7564 5636
rect 7392 5596 7564 5624
rect 7558 5584 7564 5596
rect 7616 5624 7622 5636
rect 7760 5624 7788 5655
rect 8018 5652 8024 5704
rect 8076 5692 8082 5704
rect 8481 5695 8539 5701
rect 8481 5692 8493 5695
rect 8076 5664 8493 5692
rect 8076 5652 8082 5664
rect 8481 5661 8493 5664
rect 8527 5661 8539 5695
rect 8481 5655 8539 5661
rect 7616 5596 8156 5624
rect 7616 5584 7622 5596
rect 8128 5568 8156 5596
rect 2004 5528 3188 5556
rect 4433 5559 4491 5565
rect 2004 5516 2010 5528
rect 4433 5525 4445 5559
rect 4479 5525 4491 5559
rect 4433 5519 4491 5525
rect 4522 5516 4528 5568
rect 4580 5556 4586 5568
rect 4801 5559 4859 5565
rect 4801 5556 4813 5559
rect 4580 5528 4813 5556
rect 4580 5516 4586 5528
rect 4801 5525 4813 5528
rect 4847 5525 4859 5559
rect 4801 5519 4859 5525
rect 8110 5516 8116 5568
rect 8168 5516 8174 5568
rect 1104 5466 9384 5488
rect 1104 5414 2645 5466
rect 2697 5414 2709 5466
rect 2761 5414 2773 5466
rect 2825 5414 2837 5466
rect 2889 5414 2901 5466
rect 2953 5414 4715 5466
rect 4767 5414 4779 5466
rect 4831 5414 4843 5466
rect 4895 5414 4907 5466
rect 4959 5414 4971 5466
rect 5023 5414 6785 5466
rect 6837 5414 6849 5466
rect 6901 5414 6913 5466
rect 6965 5414 6977 5466
rect 7029 5414 7041 5466
rect 7093 5414 8855 5466
rect 8907 5414 8919 5466
rect 8971 5414 8983 5466
rect 9035 5414 9047 5466
rect 9099 5414 9111 5466
rect 9163 5414 9384 5466
rect 1104 5392 9384 5414
rect 1394 5312 1400 5364
rect 1452 5312 1458 5364
rect 1762 5312 1768 5364
rect 1820 5312 1826 5364
rect 2314 5312 2320 5364
rect 2372 5312 2378 5364
rect 5074 5312 5080 5364
rect 5132 5312 5138 5364
rect 8018 5312 8024 5364
rect 8076 5312 8082 5364
rect 1412 5284 1440 5312
rect 1673 5287 1731 5293
rect 1673 5284 1685 5287
rect 1412 5256 1685 5284
rect 1673 5253 1685 5256
rect 1719 5253 1731 5287
rect 2332 5284 2360 5312
rect 2685 5287 2743 5293
rect 2685 5284 2697 5287
rect 1673 5247 1731 5253
rect 1872 5256 2176 5284
rect 2332 5256 2697 5284
rect 1397 5219 1455 5225
rect 1397 5185 1409 5219
rect 1443 5185 1455 5219
rect 1397 5179 1455 5185
rect 1489 5219 1547 5225
rect 1489 5185 1501 5219
rect 1535 5216 1547 5219
rect 1578 5216 1584 5228
rect 1535 5188 1584 5216
rect 1535 5185 1547 5188
rect 1489 5179 1547 5185
rect 1412 5148 1440 5179
rect 1578 5176 1584 5188
rect 1636 5216 1642 5228
rect 1872 5216 1900 5256
rect 1636 5188 1900 5216
rect 1636 5176 1642 5188
rect 1946 5176 1952 5228
rect 2004 5176 2010 5228
rect 2041 5219 2099 5225
rect 2041 5185 2053 5219
rect 2087 5185 2099 5219
rect 2148 5216 2176 5256
rect 2685 5253 2697 5256
rect 2731 5253 2743 5287
rect 5092 5284 5120 5312
rect 2685 5247 2743 5253
rect 4448 5256 4752 5284
rect 5092 5256 5488 5284
rect 4448 5228 4476 5256
rect 2317 5219 2375 5225
rect 2317 5216 2329 5219
rect 2148 5188 2329 5216
rect 2041 5179 2099 5185
rect 2317 5185 2329 5188
rect 2363 5185 2375 5219
rect 2317 5179 2375 5185
rect 2056 5148 2084 5179
rect 2866 5176 2872 5228
rect 2924 5176 2930 5228
rect 4430 5176 4436 5228
rect 4488 5176 4494 5228
rect 4617 5219 4675 5225
rect 4617 5185 4629 5219
rect 4663 5185 4675 5219
rect 4724 5216 4752 5256
rect 5077 5219 5135 5225
rect 5077 5216 5089 5219
rect 4724 5188 5089 5216
rect 4617 5179 4675 5185
rect 5077 5185 5089 5188
rect 5123 5185 5135 5219
rect 5077 5179 5135 5185
rect 5261 5219 5319 5225
rect 5261 5185 5273 5219
rect 5307 5185 5319 5219
rect 5261 5179 5319 5185
rect 1412 5120 1532 5148
rect 1504 5012 1532 5120
rect 1688 5120 2084 5148
rect 1688 5089 1716 5120
rect 2130 5108 2136 5160
rect 2188 5108 2194 5160
rect 4522 5108 4528 5160
rect 4580 5108 4586 5160
rect 4632 5148 4660 5179
rect 5276 5148 5304 5179
rect 5350 5176 5356 5228
rect 5408 5176 5414 5228
rect 5460 5225 5488 5256
rect 5445 5219 5503 5225
rect 5445 5185 5457 5219
rect 5491 5185 5503 5219
rect 5445 5179 5503 5185
rect 5626 5176 5632 5228
rect 5684 5216 5690 5228
rect 7653 5219 7711 5225
rect 7653 5216 7665 5219
rect 5684 5188 7665 5216
rect 5684 5176 5690 5188
rect 7653 5185 7665 5188
rect 7699 5216 7711 5219
rect 7699 5188 8064 5216
rect 7699 5185 7711 5188
rect 7653 5179 7711 5185
rect 8036 5160 8064 5188
rect 8202 5176 8208 5228
rect 8260 5216 8266 5228
rect 8757 5219 8815 5225
rect 8757 5216 8769 5219
rect 8260 5188 8769 5216
rect 8260 5176 8266 5188
rect 8757 5185 8769 5188
rect 8803 5185 8815 5219
rect 8757 5179 8815 5185
rect 4632 5120 5488 5148
rect 1673 5083 1731 5089
rect 1673 5049 1685 5083
rect 1719 5049 1731 5083
rect 1673 5043 1731 5049
rect 2148 5080 2176 5108
rect 2225 5083 2283 5089
rect 2225 5080 2237 5083
rect 2148 5052 2237 5080
rect 2148 5012 2176 5052
rect 2225 5049 2237 5052
rect 2271 5049 2283 5083
rect 2225 5043 2283 5049
rect 3418 5040 3424 5092
rect 3476 5080 3482 5092
rect 4062 5080 4068 5092
rect 3476 5052 4068 5080
rect 3476 5040 3482 5052
rect 4062 5040 4068 5052
rect 4120 5080 4126 5092
rect 5166 5080 5172 5092
rect 4120 5052 5172 5080
rect 4120 5040 4126 5052
rect 5166 5040 5172 5052
rect 5224 5040 5230 5092
rect 5460 5024 5488 5120
rect 7558 5108 7564 5160
rect 7616 5108 7622 5160
rect 7742 5108 7748 5160
rect 7800 5108 7806 5160
rect 7834 5108 7840 5160
rect 7892 5108 7898 5160
rect 8018 5108 8024 5160
rect 8076 5108 8082 5160
rect 9030 5108 9036 5160
rect 9088 5108 9094 5160
rect 1504 4984 2176 5012
rect 3050 4972 3056 5024
rect 3108 4972 3114 5024
rect 4890 4972 4896 5024
rect 4948 4972 4954 5024
rect 5442 4972 5448 5024
rect 5500 4972 5506 5024
rect 5721 5015 5779 5021
rect 5721 4981 5733 5015
rect 5767 5012 5779 5015
rect 6546 5012 6552 5024
rect 5767 4984 6552 5012
rect 5767 4981 5779 4984
rect 5721 4975 5779 4981
rect 6546 4972 6552 4984
rect 6604 5012 6610 5024
rect 7190 5012 7196 5024
rect 6604 4984 7196 5012
rect 6604 4972 6610 4984
rect 7190 4972 7196 4984
rect 7248 4972 7254 5024
rect 1104 4922 9384 4944
rect 1104 4870 1985 4922
rect 2037 4870 2049 4922
rect 2101 4870 2113 4922
rect 2165 4870 2177 4922
rect 2229 4870 2241 4922
rect 2293 4870 4055 4922
rect 4107 4870 4119 4922
rect 4171 4870 4183 4922
rect 4235 4870 4247 4922
rect 4299 4870 4311 4922
rect 4363 4870 6125 4922
rect 6177 4870 6189 4922
rect 6241 4870 6253 4922
rect 6305 4870 6317 4922
rect 6369 4870 6381 4922
rect 6433 4870 8195 4922
rect 8247 4870 8259 4922
rect 8311 4870 8323 4922
rect 8375 4870 8387 4922
rect 8439 4870 8451 4922
rect 8503 4870 9384 4922
rect 1104 4848 9384 4870
rect 2593 4811 2651 4817
rect 2593 4777 2605 4811
rect 2639 4808 2651 4811
rect 2866 4808 2872 4820
rect 2639 4780 2872 4808
rect 2639 4777 2651 4780
rect 2593 4771 2651 4777
rect 2866 4768 2872 4780
rect 2924 4768 2930 4820
rect 4890 4768 4896 4820
rect 4948 4768 4954 4820
rect 5442 4768 5448 4820
rect 5500 4768 5506 4820
rect 7098 4808 7104 4820
rect 6748 4780 7104 4808
rect 1673 4743 1731 4749
rect 1673 4709 1685 4743
rect 1719 4740 1731 4743
rect 2958 4740 2964 4752
rect 1719 4712 2964 4740
rect 1719 4709 1731 4712
rect 1673 4703 1731 4709
rect 2958 4700 2964 4712
rect 3016 4700 3022 4752
rect 2590 4632 2596 4684
rect 2648 4672 2654 4684
rect 4801 4675 4859 4681
rect 4801 4672 4813 4675
rect 2648 4644 4813 4672
rect 2648 4632 2654 4644
rect 4801 4641 4813 4644
rect 4847 4641 4859 4675
rect 4908 4672 4936 4768
rect 5534 4700 5540 4752
rect 5592 4740 5598 4752
rect 6748 4749 6776 4780
rect 7098 4768 7104 4780
rect 7156 4768 7162 4820
rect 7190 4768 7196 4820
rect 7248 4768 7254 4820
rect 7561 4811 7619 4817
rect 7561 4777 7573 4811
rect 7607 4808 7619 4811
rect 7834 4808 7840 4820
rect 7607 4780 7840 4808
rect 7607 4777 7619 4780
rect 7561 4771 7619 4777
rect 7834 4768 7840 4780
rect 7892 4768 7898 4820
rect 6733 4743 6791 4749
rect 6733 4740 6745 4743
rect 5592 4712 6745 4740
rect 5592 4700 5598 4712
rect 5629 4675 5687 4681
rect 4908 4644 5304 4672
rect 4801 4635 4859 4641
rect 934 4564 940 4616
rect 992 4604 998 4616
rect 1489 4607 1547 4613
rect 1489 4604 1501 4607
rect 992 4576 1501 4604
rect 992 4564 998 4576
rect 1489 4573 1501 4576
rect 1535 4573 1547 4607
rect 1489 4567 1547 4573
rect 1578 4564 1584 4616
rect 1636 4604 1642 4616
rect 2501 4607 2559 4613
rect 2501 4604 2513 4607
rect 1636 4576 2513 4604
rect 1636 4564 1642 4576
rect 2501 4573 2513 4576
rect 2547 4573 2559 4607
rect 2501 4567 2559 4573
rect 3050 4564 3056 4616
rect 3108 4604 3114 4616
rect 3789 4607 3847 4613
rect 3789 4604 3801 4607
rect 3108 4576 3801 4604
rect 3108 4564 3114 4576
rect 3789 4573 3801 4576
rect 3835 4573 3847 4607
rect 3789 4567 3847 4573
rect 3804 4536 3832 4567
rect 3878 4564 3884 4616
rect 3936 4604 3942 4616
rect 3973 4607 4031 4613
rect 3973 4604 3985 4607
rect 3936 4576 3985 4604
rect 3936 4564 3942 4576
rect 3973 4573 3985 4576
rect 4019 4573 4031 4607
rect 3973 4567 4031 4573
rect 4062 4564 4068 4616
rect 4120 4564 4126 4616
rect 4249 4607 4307 4613
rect 4249 4573 4261 4607
rect 4295 4573 4307 4607
rect 4249 4567 4307 4573
rect 4985 4607 5043 4613
rect 4985 4573 4997 4607
rect 5031 4604 5043 4607
rect 5074 4604 5080 4616
rect 5031 4576 5080 4604
rect 5031 4573 5043 4576
rect 4985 4567 5043 4573
rect 4264 4536 4292 4567
rect 5074 4564 5080 4576
rect 5132 4564 5138 4616
rect 5276 4613 5304 4644
rect 5629 4641 5641 4675
rect 5675 4641 5687 4675
rect 5629 4635 5687 4641
rect 5261 4607 5319 4613
rect 5261 4573 5273 4607
rect 5307 4573 5319 4607
rect 5261 4567 5319 4573
rect 5350 4536 5356 4548
rect 3804 4508 4292 4536
rect 5092 4508 5356 4536
rect 3786 4428 3792 4480
rect 3844 4428 3850 4480
rect 4249 4471 4307 4477
rect 4249 4437 4261 4471
rect 4295 4468 4307 4471
rect 5092 4468 5120 4508
rect 5350 4496 5356 4508
rect 5408 4496 5414 4548
rect 5644 4536 5672 4635
rect 5736 4613 5764 4712
rect 6733 4709 6745 4712
rect 6779 4709 6791 4743
rect 7650 4740 7656 4752
rect 6733 4703 6791 4709
rect 6840 4712 7656 4740
rect 6840 4672 6868 4712
rect 7650 4700 7656 4712
rect 7708 4740 7714 4752
rect 7708 4712 7972 4740
rect 7708 4700 7714 4712
rect 6656 4644 6868 4672
rect 6917 4675 6975 4681
rect 6656 4616 6684 4644
rect 6917 4641 6929 4675
rect 6963 4672 6975 4675
rect 7282 4672 7288 4684
rect 6963 4644 7288 4672
rect 6963 4641 6975 4644
rect 6917 4635 6975 4641
rect 7282 4632 7288 4644
rect 7340 4632 7346 4684
rect 5721 4607 5779 4613
rect 5721 4573 5733 4607
rect 5767 4573 5779 4607
rect 5721 4567 5779 4573
rect 6638 4564 6644 4616
rect 6696 4564 6702 4616
rect 7944 4613 7972 4712
rect 8018 4700 8024 4752
rect 8076 4740 8082 4752
rect 8205 4743 8263 4749
rect 8205 4740 8217 4743
rect 8076 4712 8217 4740
rect 8076 4700 8082 4712
rect 8205 4709 8217 4712
rect 8251 4709 8263 4743
rect 8205 4703 8263 4709
rect 7193 4607 7251 4613
rect 7193 4573 7205 4607
rect 7239 4573 7251 4607
rect 7193 4567 7251 4573
rect 7929 4607 7987 4613
rect 7929 4573 7941 4607
rect 7975 4573 7987 4607
rect 7929 4567 7987 4573
rect 6457 4539 6515 4545
rect 6457 4536 6469 4539
rect 5644 4508 6469 4536
rect 5736 4480 5764 4508
rect 6457 4505 6469 4508
rect 6503 4505 6515 4539
rect 6457 4499 6515 4505
rect 7208 4480 7236 4567
rect 8110 4564 8116 4616
rect 8168 4564 8174 4616
rect 4295 4440 5120 4468
rect 4295 4437 4307 4440
rect 4249 4431 4307 4437
rect 5166 4428 5172 4480
rect 5224 4468 5230 4480
rect 5626 4468 5632 4480
rect 5224 4440 5632 4468
rect 5224 4428 5230 4440
rect 5626 4428 5632 4440
rect 5684 4428 5690 4480
rect 5718 4428 5724 4480
rect 5776 4428 5782 4480
rect 7190 4428 7196 4480
rect 7248 4428 7254 4480
rect 1104 4378 9384 4400
rect 1104 4326 2645 4378
rect 2697 4326 2709 4378
rect 2761 4326 2773 4378
rect 2825 4326 2837 4378
rect 2889 4326 2901 4378
rect 2953 4326 4715 4378
rect 4767 4326 4779 4378
rect 4831 4326 4843 4378
rect 4895 4326 4907 4378
rect 4959 4326 4971 4378
rect 5023 4326 6785 4378
rect 6837 4326 6849 4378
rect 6901 4326 6913 4378
rect 6965 4326 6977 4378
rect 7029 4326 7041 4378
rect 7093 4326 8855 4378
rect 8907 4326 8919 4378
rect 8971 4326 8983 4378
rect 9035 4326 9047 4378
rect 9099 4326 9111 4378
rect 9163 4326 9384 4378
rect 1104 4304 9384 4326
rect 3252 4236 3556 4264
rect 1670 4088 1676 4140
rect 1728 4088 1734 4140
rect 1854 4088 1860 4140
rect 1912 4088 1918 4140
rect 2041 4131 2099 4137
rect 2041 4097 2053 4131
rect 2087 4097 2099 4131
rect 2041 4091 2099 4097
rect 2133 4131 2191 4137
rect 2133 4097 2145 4131
rect 2179 4097 2191 4131
rect 2133 4091 2191 4097
rect 2869 4131 2927 4137
rect 2869 4097 2881 4131
rect 2915 4097 2927 4131
rect 2869 4091 2927 4097
rect 3053 4131 3111 4137
rect 3053 4097 3065 4131
rect 3099 4128 3111 4131
rect 3252 4128 3280 4236
rect 3099 4100 3280 4128
rect 3329 4131 3387 4137
rect 3099 4097 3111 4100
rect 3053 4091 3111 4097
rect 3329 4097 3341 4131
rect 3375 4126 3387 4131
rect 3418 4126 3424 4140
rect 3375 4098 3424 4126
rect 3375 4097 3387 4098
rect 3329 4091 3387 4097
rect 2056 3924 2084 4091
rect 2148 3992 2176 4091
rect 2884 4060 2912 4091
rect 3418 4088 3424 4098
rect 3476 4088 3482 4140
rect 3528 4137 3556 4236
rect 7282 4224 7288 4276
rect 7340 4224 7346 4276
rect 3513 4131 3571 4137
rect 3513 4097 3525 4131
rect 3559 4128 3571 4131
rect 3786 4128 3792 4140
rect 3559 4100 3792 4128
rect 3559 4097 3571 4100
rect 3513 4091 3571 4097
rect 3786 4088 3792 4100
rect 3844 4088 3850 4140
rect 3881 4131 3939 4137
rect 3881 4097 3893 4131
rect 3927 4128 3939 4131
rect 4430 4128 4436 4140
rect 3927 4100 4436 4128
rect 3927 4097 3939 4100
rect 3881 4091 3939 4097
rect 3605 4063 3663 4069
rect 3605 4060 3617 4063
rect 2884 4032 3617 4060
rect 3605 4029 3617 4032
rect 3651 4060 3663 4063
rect 3697 4063 3755 4069
rect 3697 4060 3709 4063
rect 3651 4032 3709 4060
rect 3651 4029 3663 4032
rect 3605 4023 3663 4029
rect 3697 4029 3709 4032
rect 3743 4029 3755 4063
rect 3697 4023 3755 4029
rect 3145 3995 3203 4001
rect 3145 3992 3157 3995
rect 2148 3964 3157 3992
rect 3145 3961 3157 3964
rect 3191 3961 3203 3995
rect 3896 3992 3924 4091
rect 4430 4088 4436 4100
rect 4488 4088 4494 4140
rect 6546 4088 6552 4140
rect 6604 4088 6610 4140
rect 7009 4131 7067 4137
rect 7009 4097 7021 4131
rect 7055 4128 7067 4131
rect 7300 4128 7328 4224
rect 7055 4100 7328 4128
rect 7055 4097 7067 4100
rect 7009 4091 7067 4097
rect 3970 4020 3976 4072
rect 4028 4060 4034 4072
rect 4065 4063 4123 4069
rect 4065 4060 4077 4063
rect 4028 4032 4077 4060
rect 4028 4020 4034 4032
rect 4065 4029 4077 4032
rect 4111 4029 4123 4063
rect 6564 4060 6592 4088
rect 7101 4063 7159 4069
rect 7101 4060 7113 4063
rect 6564 4032 7113 4060
rect 4065 4023 4123 4029
rect 7101 4029 7113 4032
rect 7147 4029 7159 4063
rect 7101 4023 7159 4029
rect 7282 4020 7288 4072
rect 7340 4020 7346 4072
rect 7742 4020 7748 4072
rect 7800 4020 7806 4072
rect 3145 3955 3203 3961
rect 3436 3964 3924 3992
rect 7193 3995 7251 4001
rect 3436 3936 3464 3964
rect 7193 3961 7205 3995
rect 7239 3992 7251 3995
rect 7760 3992 7788 4020
rect 7239 3964 7788 3992
rect 7239 3961 7251 3964
rect 7193 3955 7251 3961
rect 2961 3927 3019 3933
rect 2961 3924 2973 3927
rect 2056 3896 2973 3924
rect 2961 3893 2973 3896
rect 3007 3893 3019 3927
rect 2961 3887 3019 3893
rect 3418 3884 3424 3936
rect 3476 3884 3482 3936
rect 7374 3884 7380 3936
rect 7432 3924 7438 3936
rect 7742 3924 7748 3936
rect 7432 3896 7748 3924
rect 7432 3884 7438 3896
rect 7742 3884 7748 3896
rect 7800 3884 7806 3936
rect 1104 3834 9384 3856
rect 1104 3782 1985 3834
rect 2037 3782 2049 3834
rect 2101 3782 2113 3834
rect 2165 3782 2177 3834
rect 2229 3782 2241 3834
rect 2293 3782 4055 3834
rect 4107 3782 4119 3834
rect 4171 3782 4183 3834
rect 4235 3782 4247 3834
rect 4299 3782 4311 3834
rect 4363 3782 6125 3834
rect 6177 3782 6189 3834
rect 6241 3782 6253 3834
rect 6305 3782 6317 3834
rect 6369 3782 6381 3834
rect 6433 3782 8195 3834
rect 8247 3782 8259 3834
rect 8311 3782 8323 3834
rect 8375 3782 8387 3834
rect 8439 3782 8451 3834
rect 8503 3782 9384 3834
rect 1104 3760 9384 3782
rect 1578 3680 1584 3732
rect 1636 3680 1642 3732
rect 1765 3723 1823 3729
rect 1765 3689 1777 3723
rect 1811 3720 1823 3723
rect 1854 3720 1860 3732
rect 1811 3692 1860 3720
rect 1811 3689 1823 3692
rect 1765 3683 1823 3689
rect 1854 3680 1860 3692
rect 1912 3680 1918 3732
rect 3513 3723 3571 3729
rect 3513 3689 3525 3723
rect 3559 3720 3571 3723
rect 3970 3720 3976 3732
rect 3559 3692 3976 3720
rect 3559 3689 3571 3692
rect 3513 3683 3571 3689
rect 3970 3680 3976 3692
rect 4028 3680 4034 3732
rect 5074 3680 5080 3732
rect 5132 3680 5138 3732
rect 5534 3680 5540 3732
rect 5592 3680 5598 3732
rect 1964 3624 2268 3652
rect 1964 3593 1992 3624
rect 1949 3587 2007 3593
rect 1949 3553 1961 3587
rect 1995 3553 2007 3587
rect 1949 3547 2007 3553
rect 2130 3544 2136 3596
rect 2188 3544 2194 3596
rect 2240 3584 2268 3624
rect 4338 3612 4344 3664
rect 4396 3612 4402 3664
rect 2406 3584 2412 3596
rect 2240 3556 2412 3584
rect 2406 3544 2412 3556
rect 2464 3584 2470 3596
rect 5445 3587 5503 3593
rect 2464 3556 5304 3584
rect 2464 3544 2470 3556
rect 2041 3519 2099 3525
rect 2041 3485 2053 3519
rect 2087 3485 2099 3519
rect 2041 3479 2099 3485
rect 934 3408 940 3460
rect 992 3448 998 3460
rect 1489 3451 1547 3457
rect 1489 3448 1501 3451
rect 992 3420 1501 3448
rect 992 3408 998 3420
rect 1489 3417 1501 3420
rect 1535 3417 1547 3451
rect 2056 3448 2084 3479
rect 2222 3476 2228 3528
rect 2280 3476 2286 3528
rect 3234 3476 3240 3528
rect 3292 3516 3298 3528
rect 4341 3519 4399 3525
rect 4341 3516 4353 3519
rect 3292 3488 4353 3516
rect 3292 3476 3298 3488
rect 4341 3485 4353 3488
rect 4387 3516 4399 3519
rect 4430 3516 4436 3528
rect 4387 3488 4436 3516
rect 4387 3485 4399 3488
rect 4341 3479 4399 3485
rect 4430 3476 4436 3488
rect 4488 3476 4494 3528
rect 4614 3476 4620 3528
rect 4672 3476 4678 3528
rect 5276 3525 5304 3556
rect 5445 3553 5457 3587
rect 5491 3584 5503 3587
rect 5552 3584 5580 3680
rect 8481 3655 8539 3661
rect 8481 3621 8493 3655
rect 8527 3621 8539 3655
rect 8481 3615 8539 3621
rect 5491 3556 5580 3584
rect 5491 3553 5503 3556
rect 5445 3547 5503 3553
rect 7374 3544 7380 3596
rect 7432 3544 7438 3596
rect 7466 3544 7472 3596
rect 7524 3584 7530 3596
rect 7653 3587 7711 3593
rect 7653 3584 7665 3587
rect 7524 3556 7665 3584
rect 7524 3544 7530 3556
rect 7653 3553 7665 3556
rect 7699 3553 7711 3587
rect 7653 3547 7711 3553
rect 5261 3519 5319 3525
rect 5261 3485 5273 3519
rect 5307 3485 5319 3519
rect 5261 3479 5319 3485
rect 2056 3420 3096 3448
rect 1489 3411 1547 3417
rect 3068 3392 3096 3420
rect 3142 3408 3148 3460
rect 3200 3408 3206 3460
rect 3326 3408 3332 3460
rect 3384 3408 3390 3460
rect 5276 3448 5304 3479
rect 5350 3476 5356 3528
rect 5408 3476 5414 3528
rect 5534 3476 5540 3528
rect 5592 3476 5598 3528
rect 7190 3476 7196 3528
rect 7248 3516 7254 3528
rect 7745 3519 7803 3525
rect 7745 3516 7757 3519
rect 7248 3488 7757 3516
rect 7248 3476 7254 3488
rect 7745 3485 7757 3488
rect 7791 3516 7803 3519
rect 8496 3516 8524 3615
rect 7791 3488 8524 3516
rect 7791 3485 7803 3488
rect 7745 3479 7803 3485
rect 8662 3476 8668 3528
rect 8720 3476 8726 3528
rect 5276 3420 7788 3448
rect 7760 3392 7788 3420
rect 3050 3340 3056 3392
rect 3108 3380 3114 3392
rect 4525 3383 4583 3389
rect 4525 3380 4537 3383
rect 3108 3352 4537 3380
rect 3108 3340 3114 3352
rect 4525 3349 4537 3352
rect 4571 3380 4583 3383
rect 5074 3380 5080 3392
rect 4571 3352 5080 3380
rect 4571 3349 4583 3352
rect 4525 3343 4583 3349
rect 5074 3340 5080 3352
rect 5132 3340 5138 3392
rect 7742 3340 7748 3392
rect 7800 3340 7806 3392
rect 1104 3290 9384 3312
rect 1104 3238 2645 3290
rect 2697 3238 2709 3290
rect 2761 3238 2773 3290
rect 2825 3238 2837 3290
rect 2889 3238 2901 3290
rect 2953 3238 4715 3290
rect 4767 3238 4779 3290
rect 4831 3238 4843 3290
rect 4895 3238 4907 3290
rect 4959 3238 4971 3290
rect 5023 3238 6785 3290
rect 6837 3238 6849 3290
rect 6901 3238 6913 3290
rect 6965 3238 6977 3290
rect 7029 3238 7041 3290
rect 7093 3238 8855 3290
rect 8907 3238 8919 3290
rect 8971 3238 8983 3290
rect 9035 3238 9047 3290
rect 9099 3238 9111 3290
rect 9163 3238 9384 3290
rect 1104 3216 9384 3238
rect 1486 3136 1492 3188
rect 1544 3176 1550 3188
rect 1765 3179 1823 3185
rect 1765 3176 1777 3179
rect 1544 3148 1777 3176
rect 1544 3136 1550 3148
rect 1765 3145 1777 3148
rect 1811 3145 1823 3179
rect 1765 3139 1823 3145
rect 1394 3068 1400 3120
rect 1452 3108 1458 3120
rect 1581 3111 1639 3117
rect 1581 3108 1593 3111
rect 1452 3080 1593 3108
rect 1452 3068 1458 3080
rect 1581 3077 1593 3080
rect 1627 3077 1639 3111
rect 1780 3108 1808 3139
rect 2222 3136 2228 3188
rect 2280 3176 2286 3188
rect 2501 3179 2559 3185
rect 2501 3176 2513 3179
rect 2280 3148 2513 3176
rect 2280 3136 2286 3148
rect 2501 3145 2513 3148
rect 2547 3145 2559 3179
rect 2501 3139 2559 3145
rect 3142 3136 3148 3188
rect 3200 3136 3206 3188
rect 3326 3136 3332 3188
rect 3384 3136 3390 3188
rect 3418 3136 3424 3188
rect 3476 3136 3482 3188
rect 4338 3136 4344 3188
rect 4396 3136 4402 3188
rect 4430 3136 4436 3188
rect 4488 3176 4494 3188
rect 4488 3148 4936 3176
rect 4488 3136 4494 3148
rect 2130 3108 2136 3120
rect 1780 3080 2136 3108
rect 1581 3071 1639 3077
rect 1854 3000 1860 3052
rect 1912 3000 1918 3052
rect 1964 3049 1992 3080
rect 2130 3068 2136 3080
rect 2188 3068 2194 3120
rect 3050 3068 3056 3120
rect 3108 3068 3114 3120
rect 1949 3043 2007 3049
rect 1949 3009 1961 3043
rect 1995 3009 2007 3043
rect 1949 3003 2007 3009
rect 2225 3043 2283 3049
rect 2225 3009 2237 3043
rect 2271 3009 2283 3043
rect 2225 3003 2283 3009
rect 2240 2972 2268 3003
rect 2314 3000 2320 3052
rect 2372 3000 2378 3052
rect 2777 3043 2835 3049
rect 2777 3009 2789 3043
rect 2823 3040 2835 3043
rect 3068 3040 3096 3068
rect 2823 3012 3096 3040
rect 3160 3040 3188 3136
rect 3344 3108 3372 3136
rect 3605 3111 3663 3117
rect 3605 3108 3617 3111
rect 3344 3080 3617 3108
rect 3237 3043 3295 3049
rect 3237 3040 3249 3043
rect 3160 3012 3249 3040
rect 2823 3009 2835 3012
rect 2777 3003 2835 3009
rect 1596 2944 2268 2972
rect 1596 2913 1624 2944
rect 1581 2907 1639 2913
rect 1581 2873 1593 2907
rect 1627 2873 1639 2907
rect 1581 2867 1639 2873
rect 1854 2864 1860 2916
rect 1912 2904 1918 2916
rect 2041 2907 2099 2913
rect 2041 2904 2053 2907
rect 1912 2876 2053 2904
rect 1912 2864 1918 2876
rect 2041 2873 2053 2876
rect 2087 2904 2099 2907
rect 2792 2904 2820 3003
rect 2869 2975 2927 2981
rect 2869 2941 2881 2975
rect 2915 2972 2927 2975
rect 3050 2972 3056 2984
rect 2915 2944 3056 2972
rect 2915 2941 2927 2944
rect 2869 2935 2927 2941
rect 3050 2932 3056 2944
rect 3108 2932 3114 2984
rect 3160 2981 3188 3012
rect 3237 3009 3249 3012
rect 3283 3009 3295 3043
rect 3344 3040 3372 3080
rect 3605 3077 3617 3080
rect 3651 3077 3663 3111
rect 3605 3071 3663 3077
rect 3421 3043 3479 3049
rect 3421 3040 3433 3043
rect 3344 3012 3433 3040
rect 3237 3003 3295 3009
rect 3421 3009 3433 3012
rect 3467 3009 3479 3043
rect 3421 3003 3479 3009
rect 3513 3043 3571 3049
rect 3513 3009 3525 3043
rect 3559 3009 3571 3043
rect 3513 3003 3571 3009
rect 4249 3043 4307 3049
rect 4249 3009 4261 3043
rect 4295 3009 4307 3043
rect 4249 3003 4307 3009
rect 3145 2975 3203 2981
rect 3145 2941 3157 2975
rect 3191 2972 3203 2975
rect 3191 2944 3225 2972
rect 3191 2941 3203 2944
rect 3145 2935 3203 2941
rect 3528 2904 3556 3003
rect 2087 2876 2820 2904
rect 3160 2876 3556 2904
rect 4264 2904 4292 3003
rect 4356 2981 4384 3136
rect 4614 3000 4620 3052
rect 4672 3040 4678 3052
rect 4908 3049 4936 3148
rect 5534 3136 5540 3188
rect 5592 3176 5598 3188
rect 5905 3179 5963 3185
rect 5905 3176 5917 3179
rect 5592 3148 5917 3176
rect 5592 3136 5598 3148
rect 5905 3145 5917 3148
rect 5951 3145 5963 3179
rect 5905 3139 5963 3145
rect 7193 3179 7251 3185
rect 7193 3145 7205 3179
rect 7239 3176 7251 3179
rect 7282 3176 7288 3188
rect 7239 3148 7288 3176
rect 7239 3145 7251 3148
rect 7193 3139 7251 3145
rect 7282 3136 7288 3148
rect 7340 3136 7346 3188
rect 7374 3136 7380 3188
rect 7432 3136 7438 3188
rect 7558 3136 7564 3188
rect 7616 3176 7622 3188
rect 7837 3179 7895 3185
rect 7837 3176 7849 3179
rect 7616 3148 7849 3176
rect 7616 3136 7622 3148
rect 7837 3145 7849 3148
rect 7883 3145 7895 3179
rect 7837 3139 7895 3145
rect 8113 3179 8171 3185
rect 8113 3145 8125 3179
rect 8159 3176 8171 3179
rect 8570 3176 8576 3188
rect 8159 3148 8576 3176
rect 8159 3145 8171 3148
rect 8113 3139 8171 3145
rect 8570 3136 8576 3148
rect 8628 3136 8634 3188
rect 5261 3111 5319 3117
rect 5261 3077 5273 3111
rect 5307 3108 5319 3111
rect 5307 3080 6868 3108
rect 5307 3077 5319 3080
rect 5261 3071 5319 3077
rect 4801 3043 4859 3049
rect 4801 3040 4813 3043
rect 4672 3012 4813 3040
rect 4672 3000 4678 3012
rect 4801 3009 4813 3012
rect 4847 3009 4859 3043
rect 4801 3003 4859 3009
rect 4893 3043 4951 3049
rect 4893 3009 4905 3043
rect 4939 3009 4951 3043
rect 4893 3003 4951 3009
rect 5074 3000 5080 3052
rect 5132 3000 5138 3052
rect 5353 3043 5411 3049
rect 5353 3009 5365 3043
rect 5399 3040 5411 3043
rect 5442 3040 5448 3052
rect 5399 3012 5448 3040
rect 5399 3009 5411 3012
rect 5353 3003 5411 3009
rect 5442 3000 5448 3012
rect 5500 3000 5506 3052
rect 5626 3000 5632 3052
rect 5684 3000 5690 3052
rect 5721 3043 5779 3049
rect 5721 3009 5733 3043
rect 5767 3040 5779 3043
rect 6454 3040 6460 3052
rect 5767 3012 6460 3040
rect 5767 3009 5779 3012
rect 5721 3003 5779 3009
rect 6454 3000 6460 3012
rect 6512 3000 6518 3052
rect 6840 3049 6868 3080
rect 6825 3043 6883 3049
rect 6825 3009 6837 3043
rect 6871 3009 6883 3043
rect 6825 3003 6883 3009
rect 7190 3000 7196 3052
rect 7248 3040 7254 3052
rect 7285 3043 7343 3049
rect 7285 3040 7297 3043
rect 7248 3012 7297 3040
rect 7248 3000 7254 3012
rect 7285 3009 7297 3012
rect 7331 3009 7343 3043
rect 7285 3003 7343 3009
rect 4341 2975 4399 2981
rect 4341 2941 4353 2975
rect 4387 2941 4399 2975
rect 4341 2935 4399 2941
rect 4430 2932 4436 2984
rect 4488 2972 4494 2984
rect 5092 2972 5120 3000
rect 4488 2944 5028 2972
rect 5092 2944 5856 2972
rect 4488 2932 4494 2944
rect 4448 2904 4476 2932
rect 5000 2913 5028 2944
rect 4264 2876 4476 2904
rect 4985 2907 5043 2913
rect 2087 2873 2099 2876
rect 2041 2867 2099 2873
rect 2130 2796 2136 2848
rect 2188 2836 2194 2848
rect 3160 2836 3188 2876
rect 4985 2873 4997 2907
rect 5031 2904 5043 2907
rect 5350 2904 5356 2916
rect 5031 2876 5356 2904
rect 5031 2873 5043 2876
rect 4985 2867 5043 2873
rect 5350 2864 5356 2876
rect 5408 2904 5414 2916
rect 5445 2907 5503 2913
rect 5445 2904 5457 2907
rect 5408 2876 5457 2904
rect 5408 2864 5414 2876
rect 5445 2873 5457 2876
rect 5491 2873 5503 2907
rect 5445 2867 5503 2873
rect 2188 2808 3188 2836
rect 4525 2839 4583 2845
rect 2188 2796 2194 2808
rect 4525 2805 4537 2839
rect 4571 2836 4583 2839
rect 5718 2836 5724 2848
rect 4571 2808 5724 2836
rect 4571 2805 4583 2808
rect 4525 2799 4583 2805
rect 5718 2796 5724 2808
rect 5776 2796 5782 2848
rect 5828 2836 5856 2944
rect 6472 2904 6500 3000
rect 6917 2975 6975 2981
rect 6917 2941 6929 2975
rect 6963 2972 6975 2975
rect 7392 2972 7420 3136
rect 7558 3000 7564 3052
rect 7616 3000 7622 3052
rect 7653 3043 7711 3049
rect 7653 3009 7665 3043
rect 7699 3009 7711 3043
rect 7653 3003 7711 3009
rect 6963 2944 7420 2972
rect 6963 2941 6975 2944
rect 6917 2935 6975 2941
rect 7668 2904 7696 3003
rect 7926 3000 7932 3052
rect 7984 3000 7990 3052
rect 8110 3000 8116 3052
rect 8168 3040 8174 3052
rect 8757 3043 8815 3049
rect 8757 3040 8769 3043
rect 8168 3012 8769 3040
rect 8168 3000 8174 3012
rect 8757 3009 8769 3012
rect 8803 3009 8815 3043
rect 8757 3003 8815 3009
rect 8941 3043 8999 3049
rect 8941 3009 8953 3043
rect 8987 3040 8999 3043
rect 9398 3040 9404 3052
rect 8987 3012 9404 3040
rect 8987 3009 8999 3012
rect 8941 3003 8999 3009
rect 9398 3000 9404 3012
rect 9456 3000 9462 3052
rect 6472 2876 7696 2904
rect 6730 2836 6736 2848
rect 5828 2808 6736 2836
rect 6730 2796 6736 2808
rect 6788 2796 6794 2848
rect 7374 2796 7380 2848
rect 7432 2796 7438 2848
rect 1104 2746 9384 2768
rect 1104 2694 1985 2746
rect 2037 2694 2049 2746
rect 2101 2694 2113 2746
rect 2165 2694 2177 2746
rect 2229 2694 2241 2746
rect 2293 2694 4055 2746
rect 4107 2694 4119 2746
rect 4171 2694 4183 2746
rect 4235 2694 4247 2746
rect 4299 2694 4311 2746
rect 4363 2694 6125 2746
rect 6177 2694 6189 2746
rect 6241 2694 6253 2746
rect 6305 2694 6317 2746
rect 6369 2694 6381 2746
rect 6433 2694 8195 2746
rect 8247 2694 8259 2746
rect 8311 2694 8323 2746
rect 8375 2694 8387 2746
rect 8439 2694 8451 2746
rect 8503 2694 9384 2746
rect 1104 2672 9384 2694
rect 2501 2635 2559 2641
rect 2501 2601 2513 2635
rect 2547 2632 2559 2635
rect 3510 2632 3516 2644
rect 2547 2604 3516 2632
rect 2547 2601 2559 2604
rect 2501 2595 2559 2601
rect 3510 2592 3516 2604
rect 3568 2592 3574 2644
rect 4430 2632 4436 2644
rect 3988 2604 4436 2632
rect 1673 2567 1731 2573
rect 1673 2533 1685 2567
rect 1719 2564 1731 2567
rect 3988 2564 4016 2604
rect 4430 2592 4436 2604
rect 4488 2592 4494 2644
rect 5626 2592 5632 2644
rect 5684 2632 5690 2644
rect 5721 2635 5779 2641
rect 5721 2632 5733 2635
rect 5684 2604 5733 2632
rect 5684 2592 5690 2604
rect 5721 2601 5733 2604
rect 5767 2601 5779 2635
rect 5721 2595 5779 2601
rect 5994 2592 6000 2644
rect 6052 2592 6058 2644
rect 6638 2592 6644 2644
rect 6696 2592 6702 2644
rect 7377 2635 7435 2641
rect 7377 2601 7389 2635
rect 7423 2632 7435 2635
rect 7558 2632 7564 2644
rect 7423 2604 7564 2632
rect 7423 2601 7435 2604
rect 7377 2595 7435 2601
rect 7558 2592 7564 2604
rect 7616 2592 7622 2644
rect 8573 2635 8631 2641
rect 8573 2632 8585 2635
rect 7668 2604 8585 2632
rect 1719 2536 4016 2564
rect 4065 2567 4123 2573
rect 1719 2533 1731 2536
rect 1673 2527 1731 2533
rect 4065 2533 4077 2567
rect 4111 2564 4123 2567
rect 6656 2564 6684 2592
rect 4111 2536 6684 2564
rect 4111 2533 4123 2536
rect 4065 2527 4123 2533
rect 6730 2524 6736 2576
rect 6788 2564 6794 2576
rect 7668 2564 7696 2604
rect 8573 2601 8585 2604
rect 8619 2601 8631 2635
rect 8573 2595 8631 2601
rect 6788 2536 7696 2564
rect 8021 2567 8079 2573
rect 6788 2524 6794 2536
rect 8021 2533 8033 2567
rect 8067 2533 8079 2567
rect 8021 2527 8079 2533
rect 1302 2456 1308 2508
rect 1360 2496 1366 2508
rect 2961 2499 3019 2505
rect 1360 2468 2728 2496
rect 1360 2456 1366 2468
rect 1210 2388 1216 2440
rect 1268 2428 1274 2440
rect 2700 2437 2728 2468
rect 2961 2465 2973 2499
rect 3007 2496 3019 2499
rect 3007 2468 6914 2496
rect 3007 2465 3019 2468
rect 2961 2459 3019 2465
rect 2317 2431 2375 2437
rect 2317 2428 2329 2431
rect 1268 2400 2329 2428
rect 1268 2388 1274 2400
rect 2317 2397 2329 2400
rect 2363 2397 2375 2431
rect 2317 2391 2375 2397
rect 2685 2431 2743 2437
rect 2685 2397 2697 2431
rect 2731 2397 2743 2431
rect 2685 2391 2743 2397
rect 5442 2388 5448 2440
rect 5500 2388 5506 2440
rect 5534 2388 5540 2440
rect 5592 2388 5598 2440
rect 5810 2388 5816 2440
rect 5868 2428 5874 2440
rect 6641 2431 6699 2437
rect 6641 2428 6653 2431
rect 5868 2400 6653 2428
rect 5868 2388 5874 2400
rect 6641 2397 6653 2400
rect 6687 2397 6699 2431
rect 6641 2391 6699 2397
rect 14 2320 20 2372
rect 72 2360 78 2372
rect 1489 2363 1547 2369
rect 1489 2360 1501 2363
rect 72 2332 1501 2360
rect 72 2320 78 2332
rect 1489 2329 1501 2332
rect 1535 2329 1547 2363
rect 1489 2323 1547 2329
rect 3234 2320 3240 2372
rect 3292 2360 3298 2372
rect 3881 2363 3939 2369
rect 3881 2360 3893 2363
rect 3292 2332 3893 2360
rect 3292 2320 3298 2332
rect 3881 2329 3893 2332
rect 3927 2329 3939 2363
rect 3881 2323 3939 2329
rect 5718 2320 5724 2372
rect 5776 2320 5782 2372
rect 5905 2363 5963 2369
rect 5905 2329 5917 2363
rect 5951 2329 5963 2363
rect 6886 2360 6914 2468
rect 7190 2456 7196 2508
rect 7248 2496 7254 2508
rect 7745 2499 7803 2505
rect 7745 2496 7757 2499
rect 7248 2468 7757 2496
rect 7248 2456 7254 2468
rect 7745 2465 7757 2468
rect 7791 2465 7803 2499
rect 7745 2459 7803 2465
rect 7837 2499 7895 2505
rect 7837 2465 7849 2499
rect 7883 2496 7895 2499
rect 8036 2496 8064 2527
rect 7883 2468 8064 2496
rect 7883 2465 7895 2468
rect 7837 2459 7895 2465
rect 7558 2388 7564 2440
rect 7616 2388 7622 2440
rect 7653 2431 7711 2437
rect 7653 2397 7665 2431
rect 7699 2397 7711 2431
rect 7760 2428 7788 2459
rect 8205 2431 8263 2437
rect 8205 2428 8217 2431
rect 7760 2400 8217 2428
rect 7653 2391 7711 2397
rect 8205 2397 8217 2400
rect 8251 2397 8263 2431
rect 8205 2391 8263 2397
rect 8297 2431 8355 2437
rect 8297 2397 8309 2431
rect 8343 2397 8355 2431
rect 8297 2391 8355 2397
rect 7374 2360 7380 2372
rect 6886 2332 7380 2360
rect 5905 2323 5963 2329
rect 5626 2252 5632 2304
rect 5684 2292 5690 2304
rect 5920 2292 5948 2323
rect 7374 2320 7380 2332
rect 7432 2360 7438 2372
rect 7668 2360 7696 2391
rect 7432 2332 7696 2360
rect 7432 2320 7438 2332
rect 5684 2264 5948 2292
rect 5684 2252 5690 2264
rect 6546 2252 6552 2304
rect 6604 2292 6610 2304
rect 6917 2295 6975 2301
rect 6917 2292 6929 2295
rect 6604 2264 6929 2292
rect 6604 2252 6610 2264
rect 6917 2261 6929 2264
rect 6963 2261 6975 2295
rect 7668 2292 7696 2332
rect 7742 2320 7748 2372
rect 7800 2360 7806 2372
rect 7926 2360 7932 2372
rect 7800 2332 7932 2360
rect 7800 2320 7806 2332
rect 7926 2320 7932 2332
rect 7984 2360 7990 2372
rect 8021 2363 8079 2369
rect 8021 2360 8033 2363
rect 7984 2332 8033 2360
rect 7984 2320 7990 2332
rect 8021 2329 8033 2332
rect 8067 2329 8079 2363
rect 8021 2323 8079 2329
rect 8312 2292 8340 2391
rect 8665 2363 8723 2369
rect 8665 2329 8677 2363
rect 8711 2360 8723 2363
rect 10318 2360 10324 2372
rect 8711 2332 10324 2360
rect 8711 2329 8723 2332
rect 8665 2323 8723 2329
rect 10318 2320 10324 2332
rect 10376 2320 10382 2372
rect 7668 2264 8340 2292
rect 6917 2255 6975 2261
rect 1104 2202 9384 2224
rect 1104 2150 2645 2202
rect 2697 2150 2709 2202
rect 2761 2150 2773 2202
rect 2825 2150 2837 2202
rect 2889 2150 2901 2202
rect 2953 2150 4715 2202
rect 4767 2150 4779 2202
rect 4831 2150 4843 2202
rect 4895 2150 4907 2202
rect 4959 2150 4971 2202
rect 5023 2150 6785 2202
rect 6837 2150 6849 2202
rect 6901 2150 6913 2202
rect 6965 2150 6977 2202
rect 7029 2150 7041 2202
rect 7093 2150 8855 2202
rect 8907 2150 8919 2202
rect 8971 2150 8983 2202
rect 9035 2150 9047 2202
rect 9099 2150 9111 2202
rect 9163 2150 9384 2202
rect 1104 2128 9384 2150
rect 5718 2048 5724 2100
rect 5776 2088 5782 2100
rect 7742 2088 7748 2100
rect 5776 2060 7748 2088
rect 5776 2048 5782 2060
rect 7742 2048 7748 2060
rect 7800 2048 7806 2100
<< via1 >>
rect 1985 10310 2037 10362
rect 2049 10310 2101 10362
rect 2113 10310 2165 10362
rect 2177 10310 2229 10362
rect 2241 10310 2293 10362
rect 4055 10310 4107 10362
rect 4119 10310 4171 10362
rect 4183 10310 4235 10362
rect 4247 10310 4299 10362
rect 4311 10310 4363 10362
rect 6125 10310 6177 10362
rect 6189 10310 6241 10362
rect 6253 10310 6305 10362
rect 6317 10310 6369 10362
rect 6381 10310 6433 10362
rect 8195 10310 8247 10362
rect 8259 10310 8311 10362
rect 8323 10310 8375 10362
rect 8387 10310 8439 10362
rect 8451 10310 8503 10362
rect 4620 10208 4672 10260
rect 6736 10251 6788 10260
rect 6736 10217 6745 10251
rect 6745 10217 6779 10251
rect 6779 10217 6788 10251
rect 6736 10208 6788 10217
rect 2780 10140 2832 10192
rect 1308 10004 1360 10056
rect 2596 10004 2648 10056
rect 4160 10004 4212 10056
rect 7748 10004 7800 10056
rect 8484 10004 8536 10056
rect 8668 10004 8720 10056
rect 9680 10004 9732 10056
rect 1676 9979 1728 9988
rect 1676 9945 1685 9979
rect 1685 9945 1719 9979
rect 1719 9945 1728 9979
rect 1676 9936 1728 9945
rect 2504 9936 2556 9988
rect 5080 9936 5132 9988
rect 7288 9936 7340 9988
rect 6644 9868 6696 9920
rect 7932 9911 7984 9920
rect 7932 9877 7941 9911
rect 7941 9877 7975 9911
rect 7975 9877 7984 9911
rect 7932 9868 7984 9877
rect 8392 9911 8444 9920
rect 8392 9877 8401 9911
rect 8401 9877 8435 9911
rect 8435 9877 8444 9911
rect 8392 9868 8444 9877
rect 8760 9911 8812 9920
rect 8760 9877 8769 9911
rect 8769 9877 8803 9911
rect 8803 9877 8812 9911
rect 8760 9868 8812 9877
rect 2645 9766 2697 9818
rect 2709 9766 2761 9818
rect 2773 9766 2825 9818
rect 2837 9766 2889 9818
rect 2901 9766 2953 9818
rect 4715 9766 4767 9818
rect 4779 9766 4831 9818
rect 4843 9766 4895 9818
rect 4907 9766 4959 9818
rect 4971 9766 5023 9818
rect 6785 9766 6837 9818
rect 6849 9766 6901 9818
rect 6913 9766 6965 9818
rect 6977 9766 7029 9818
rect 7041 9766 7093 9818
rect 8855 9766 8907 9818
rect 8919 9766 8971 9818
rect 8983 9766 9035 9818
rect 9047 9766 9099 9818
rect 9111 9766 9163 9818
rect 1400 9571 1452 9580
rect 1400 9537 1409 9571
rect 1409 9537 1443 9571
rect 1443 9537 1452 9571
rect 1400 9528 1452 9537
rect 2320 9571 2372 9580
rect 2320 9537 2329 9571
rect 2329 9537 2363 9571
rect 2363 9537 2372 9571
rect 2320 9528 2372 9537
rect 1676 9503 1728 9512
rect 1676 9469 1685 9503
rect 1685 9469 1719 9503
rect 1719 9469 1728 9503
rect 1676 9460 1728 9469
rect 1768 9392 1820 9444
rect 2688 9571 2740 9580
rect 2688 9537 2697 9571
rect 2697 9537 2731 9571
rect 2731 9537 2740 9571
rect 2688 9528 2740 9537
rect 3056 9571 3108 9580
rect 3056 9537 3065 9571
rect 3065 9537 3099 9571
rect 3099 9537 3108 9571
rect 3056 9528 3108 9537
rect 3240 9528 3292 9580
rect 5080 9664 5132 9716
rect 4068 9528 4120 9580
rect 4252 9528 4304 9580
rect 8392 9664 8444 9716
rect 9404 9664 9456 9716
rect 4988 9571 5040 9580
rect 4988 9537 4997 9571
rect 4997 9537 5031 9571
rect 5031 9537 5040 9571
rect 4988 9528 5040 9537
rect 3792 9460 3844 9512
rect 3976 9460 4028 9512
rect 1400 9324 1452 9376
rect 2596 9367 2648 9376
rect 2596 9333 2605 9367
rect 2605 9333 2639 9367
rect 2639 9333 2648 9367
rect 2596 9324 2648 9333
rect 3240 9324 3292 9376
rect 4160 9392 4212 9444
rect 4620 9460 4672 9512
rect 4896 9460 4948 9512
rect 5172 9571 5224 9580
rect 5172 9537 5181 9571
rect 5181 9537 5215 9571
rect 5215 9537 5224 9571
rect 5172 9528 5224 9537
rect 5356 9571 5408 9580
rect 5356 9537 5365 9571
rect 5365 9537 5399 9571
rect 5399 9537 5408 9571
rect 5356 9528 5408 9537
rect 5724 9571 5776 9580
rect 5264 9460 5316 9512
rect 5724 9537 5734 9571
rect 5734 9537 5768 9571
rect 5768 9537 5776 9571
rect 5724 9528 5776 9537
rect 6920 9571 6972 9580
rect 6920 9537 6929 9571
rect 6929 9537 6963 9571
rect 6963 9537 6972 9571
rect 6920 9528 6972 9537
rect 7380 9571 7432 9580
rect 7380 9537 7389 9571
rect 7389 9537 7423 9571
rect 7423 9537 7432 9571
rect 7380 9528 7432 9537
rect 8760 9596 8812 9648
rect 7932 9503 7984 9512
rect 7932 9469 7941 9503
rect 7941 9469 7975 9503
rect 7975 9469 7984 9503
rect 7932 9460 7984 9469
rect 4068 9324 4120 9376
rect 5080 9324 5132 9376
rect 5816 9324 5868 9376
rect 5908 9324 5960 9376
rect 6000 9367 6052 9376
rect 6000 9333 6009 9367
rect 6009 9333 6043 9367
rect 6043 9333 6052 9367
rect 6000 9324 6052 9333
rect 7748 9324 7800 9376
rect 8116 9460 8168 9512
rect 8668 9460 8720 9512
rect 1985 9222 2037 9274
rect 2049 9222 2101 9274
rect 2113 9222 2165 9274
rect 2177 9222 2229 9274
rect 2241 9222 2293 9274
rect 4055 9222 4107 9274
rect 4119 9222 4171 9274
rect 4183 9222 4235 9274
rect 4247 9222 4299 9274
rect 4311 9222 4363 9274
rect 6125 9222 6177 9274
rect 6189 9222 6241 9274
rect 6253 9222 6305 9274
rect 6317 9222 6369 9274
rect 6381 9222 6433 9274
rect 8195 9222 8247 9274
rect 8259 9222 8311 9274
rect 8323 9222 8375 9274
rect 8387 9222 8439 9274
rect 8451 9222 8503 9274
rect 2596 9120 2648 9172
rect 2688 9120 2740 9172
rect 3240 9120 3292 9172
rect 940 8916 992 8968
rect 1768 8916 1820 8968
rect 2412 8916 2464 8968
rect 3148 9052 3200 9104
rect 3976 9052 4028 9104
rect 4712 9120 4764 9172
rect 4896 9120 4948 9172
rect 5540 9120 5592 9172
rect 5816 9163 5868 9172
rect 5816 9129 5825 9163
rect 5825 9129 5859 9163
rect 5859 9129 5868 9163
rect 5816 9120 5868 9129
rect 8576 9120 8628 9172
rect 4988 9052 5040 9104
rect 6920 9052 6972 9104
rect 7840 9052 7892 9104
rect 4160 8959 4212 8968
rect 4160 8925 4169 8959
rect 4169 8925 4203 8959
rect 4203 8925 4212 8959
rect 4160 8916 4212 8925
rect 3700 8848 3752 8900
rect 3884 8848 3936 8900
rect 5264 8916 5316 8968
rect 5448 8916 5500 8968
rect 7748 8984 7800 9036
rect 8024 9027 8076 9036
rect 8024 8993 8033 9027
rect 8033 8993 8067 9027
rect 8067 8993 8076 9027
rect 8024 8984 8076 8993
rect 6920 8916 6972 8968
rect 7932 8959 7984 8968
rect 7932 8925 7941 8959
rect 7941 8925 7975 8959
rect 7975 8925 7984 8959
rect 7932 8916 7984 8925
rect 9312 8916 9364 8968
rect 5172 8780 5224 8832
rect 6000 8780 6052 8832
rect 2645 8678 2697 8730
rect 2709 8678 2761 8730
rect 2773 8678 2825 8730
rect 2837 8678 2889 8730
rect 2901 8678 2953 8730
rect 4715 8678 4767 8730
rect 4779 8678 4831 8730
rect 4843 8678 4895 8730
rect 4907 8678 4959 8730
rect 4971 8678 5023 8730
rect 6785 8678 6837 8730
rect 6849 8678 6901 8730
rect 6913 8678 6965 8730
rect 6977 8678 7029 8730
rect 7041 8678 7093 8730
rect 8855 8678 8907 8730
rect 8919 8678 8971 8730
rect 8983 8678 9035 8730
rect 9047 8678 9099 8730
rect 9111 8678 9163 8730
rect 3700 8576 3752 8628
rect 2412 8508 2464 8560
rect 3056 8508 3108 8560
rect 3884 8508 3936 8560
rect 5172 8576 5224 8628
rect 5356 8576 5408 8628
rect 6920 8576 6972 8628
rect 7564 8576 7616 8628
rect 7932 8576 7984 8628
rect 1768 8415 1820 8424
rect 1768 8381 1777 8415
rect 1777 8381 1811 8415
rect 1811 8381 1820 8415
rect 1768 8372 1820 8381
rect 4436 8440 4488 8492
rect 5264 8440 5316 8492
rect 5356 8483 5408 8492
rect 5356 8449 5365 8483
rect 5365 8449 5399 8483
rect 5399 8449 5408 8483
rect 5356 8440 5408 8449
rect 7012 8440 7064 8492
rect 7196 8483 7248 8492
rect 7196 8449 7205 8483
rect 7205 8449 7239 8483
rect 7239 8449 7248 8483
rect 7196 8440 7248 8449
rect 3516 8372 3568 8424
rect 4528 8347 4580 8356
rect 4528 8313 4537 8347
rect 4537 8313 4571 8347
rect 4571 8313 4580 8347
rect 4528 8304 4580 8313
rect 6000 8304 6052 8356
rect 8668 8483 8720 8492
rect 8668 8449 8677 8483
rect 8677 8449 8711 8483
rect 8711 8449 8720 8483
rect 8668 8440 8720 8449
rect 8024 8372 8076 8424
rect 9036 8304 9088 8356
rect 2412 8236 2464 8288
rect 2780 8279 2832 8288
rect 2780 8245 2789 8279
rect 2789 8245 2823 8279
rect 2823 8245 2832 8279
rect 2780 8236 2832 8245
rect 3240 8236 3292 8288
rect 5908 8236 5960 8288
rect 7564 8236 7616 8288
rect 1985 8134 2037 8186
rect 2049 8134 2101 8186
rect 2113 8134 2165 8186
rect 2177 8134 2229 8186
rect 2241 8134 2293 8186
rect 4055 8134 4107 8186
rect 4119 8134 4171 8186
rect 4183 8134 4235 8186
rect 4247 8134 4299 8186
rect 4311 8134 4363 8186
rect 6125 8134 6177 8186
rect 6189 8134 6241 8186
rect 6253 8134 6305 8186
rect 6317 8134 6369 8186
rect 6381 8134 6433 8186
rect 8195 8134 8247 8186
rect 8259 8134 8311 8186
rect 8323 8134 8375 8186
rect 8387 8134 8439 8186
rect 8451 8134 8503 8186
rect 1768 8032 1820 8084
rect 5080 8075 5132 8084
rect 5080 8041 5089 8075
rect 5089 8041 5123 8075
rect 5123 8041 5132 8075
rect 5080 8032 5132 8041
rect 5448 8032 5500 8084
rect 6920 8075 6972 8084
rect 6920 8041 6929 8075
rect 6929 8041 6963 8075
rect 6963 8041 6972 8075
rect 6920 8032 6972 8041
rect 7196 8032 7248 8084
rect 7380 8032 7432 8084
rect 7564 8075 7616 8084
rect 7564 8041 7573 8075
rect 7573 8041 7607 8075
rect 7607 8041 7616 8075
rect 7564 8032 7616 8041
rect 7656 8032 7708 8084
rect 8024 8075 8076 8084
rect 8024 8041 8033 8075
rect 8033 8041 8067 8075
rect 8067 8041 8076 8075
rect 8024 8032 8076 8041
rect 8576 8032 8628 8084
rect 2780 7896 2832 7948
rect 2412 7871 2464 7880
rect 2412 7837 2421 7871
rect 2421 7837 2455 7871
rect 2455 7837 2464 7871
rect 2412 7828 2464 7837
rect 2320 7803 2372 7812
rect 2320 7769 2329 7803
rect 2329 7769 2363 7803
rect 2363 7769 2372 7803
rect 5264 7964 5316 8016
rect 4436 7896 4488 7948
rect 5448 7896 5500 7948
rect 5172 7828 5224 7880
rect 5264 7871 5316 7880
rect 5264 7837 5273 7871
rect 5273 7837 5307 7871
rect 5307 7837 5316 7871
rect 5264 7828 5316 7837
rect 5908 7896 5960 7948
rect 6000 7939 6052 7948
rect 6000 7905 6009 7939
rect 6009 7905 6043 7939
rect 6043 7905 6052 7939
rect 6000 7896 6052 7905
rect 6368 7828 6420 7880
rect 2320 7760 2372 7769
rect 6092 7760 6144 7812
rect 7196 7871 7248 7880
rect 7196 7837 7205 7871
rect 7205 7837 7239 7871
rect 7239 7837 7248 7871
rect 7196 7828 7248 7837
rect 7380 7828 7432 7880
rect 5172 7692 5224 7744
rect 5908 7692 5960 7744
rect 7012 7692 7064 7744
rect 8116 7760 8168 7812
rect 8484 7692 8536 7744
rect 2645 7590 2697 7642
rect 2709 7590 2761 7642
rect 2773 7590 2825 7642
rect 2837 7590 2889 7642
rect 2901 7590 2953 7642
rect 4715 7590 4767 7642
rect 4779 7590 4831 7642
rect 4843 7590 4895 7642
rect 4907 7590 4959 7642
rect 4971 7590 5023 7642
rect 6785 7590 6837 7642
rect 6849 7590 6901 7642
rect 6913 7590 6965 7642
rect 6977 7590 7029 7642
rect 7041 7590 7093 7642
rect 8855 7590 8907 7642
rect 8919 7590 8971 7642
rect 8983 7590 9035 7642
rect 9047 7590 9099 7642
rect 9111 7590 9163 7642
rect 2320 7488 2372 7540
rect 5356 7488 5408 7540
rect 5448 7488 5500 7540
rect 6000 7488 6052 7540
rect 8668 7488 8720 7540
rect 1768 7395 1820 7404
rect 1768 7361 1777 7395
rect 1777 7361 1811 7395
rect 1811 7361 1820 7395
rect 1768 7352 1820 7361
rect 2412 7352 2464 7404
rect 2688 7395 2740 7404
rect 2688 7361 2697 7395
rect 2697 7361 2731 7395
rect 2731 7361 2740 7395
rect 2688 7352 2740 7361
rect 3516 7352 3568 7404
rect 3240 7284 3292 7336
rect 8668 7395 8720 7404
rect 8668 7361 8677 7395
rect 8677 7361 8711 7395
rect 8711 7361 8720 7395
rect 8668 7352 8720 7361
rect 6368 7284 6420 7336
rect 7196 7284 7248 7336
rect 8576 7284 8628 7336
rect 5540 7216 5592 7268
rect 8024 7216 8076 7268
rect 8484 7259 8536 7268
rect 8484 7225 8493 7259
rect 8493 7225 8527 7259
rect 8527 7225 8536 7259
rect 8484 7216 8536 7225
rect 1492 7191 1544 7200
rect 1492 7157 1501 7191
rect 1501 7157 1535 7191
rect 1535 7157 1544 7191
rect 1492 7148 1544 7157
rect 2412 7191 2464 7200
rect 2412 7157 2421 7191
rect 2421 7157 2455 7191
rect 2455 7157 2464 7191
rect 2412 7148 2464 7157
rect 3056 7148 3108 7200
rect 5172 7148 5224 7200
rect 1985 7046 2037 7098
rect 2049 7046 2101 7098
rect 2113 7046 2165 7098
rect 2177 7046 2229 7098
rect 2241 7046 2293 7098
rect 4055 7046 4107 7098
rect 4119 7046 4171 7098
rect 4183 7046 4235 7098
rect 4247 7046 4299 7098
rect 4311 7046 4363 7098
rect 6125 7046 6177 7098
rect 6189 7046 6241 7098
rect 6253 7046 6305 7098
rect 6317 7046 6369 7098
rect 6381 7046 6433 7098
rect 8195 7046 8247 7098
rect 8259 7046 8311 7098
rect 8323 7046 8375 7098
rect 8387 7046 8439 7098
rect 8451 7046 8503 7098
rect 2136 6944 2188 6996
rect 2688 6944 2740 6996
rect 4712 6944 4764 6996
rect 6000 6944 6052 6996
rect 7380 6876 7432 6928
rect 7748 6876 7800 6928
rect 8024 6876 8076 6928
rect 2320 6808 2372 6860
rect 2412 6808 2464 6860
rect 4160 6808 4212 6860
rect 4620 6808 4672 6860
rect 1860 6740 1912 6792
rect 3884 6715 3936 6724
rect 3884 6681 3893 6715
rect 3893 6681 3927 6715
rect 3927 6681 3936 6715
rect 3884 6672 3936 6681
rect 4528 6740 4580 6792
rect 6644 6740 6696 6792
rect 7196 6740 7248 6792
rect 7656 6783 7708 6792
rect 7656 6749 7665 6783
rect 7665 6749 7699 6783
rect 7699 6749 7708 6783
rect 7656 6740 7708 6749
rect 7932 6783 7984 6792
rect 7932 6749 7941 6783
rect 7941 6749 7975 6783
rect 7975 6749 7984 6783
rect 7932 6740 7984 6749
rect 8392 6783 8444 6792
rect 8392 6749 8401 6783
rect 8401 6749 8435 6783
rect 8435 6749 8444 6783
rect 8392 6740 8444 6749
rect 3976 6604 4028 6656
rect 4344 6604 4396 6656
rect 5264 6672 5316 6724
rect 7840 6604 7892 6656
rect 8208 6647 8260 6656
rect 8208 6613 8223 6647
rect 8223 6613 8257 6647
rect 8257 6613 8260 6647
rect 8208 6604 8260 6613
rect 8484 6604 8536 6656
rect 2645 6502 2697 6554
rect 2709 6502 2761 6554
rect 2773 6502 2825 6554
rect 2837 6502 2889 6554
rect 2901 6502 2953 6554
rect 4715 6502 4767 6554
rect 4779 6502 4831 6554
rect 4843 6502 4895 6554
rect 4907 6502 4959 6554
rect 4971 6502 5023 6554
rect 6785 6502 6837 6554
rect 6849 6502 6901 6554
rect 6913 6502 6965 6554
rect 6977 6502 7029 6554
rect 7041 6502 7093 6554
rect 8855 6502 8907 6554
rect 8919 6502 8971 6554
rect 8983 6502 9035 6554
rect 9047 6502 9099 6554
rect 9111 6502 9163 6554
rect 1860 6400 1912 6452
rect 4344 6400 4396 6452
rect 2136 6332 2188 6384
rect 3240 6332 3292 6384
rect 2412 6307 2464 6316
rect 2412 6273 2421 6307
rect 2421 6273 2455 6307
rect 2455 6273 2464 6307
rect 2412 6264 2464 6273
rect 3976 6332 4028 6384
rect 4160 6264 4212 6316
rect 6000 6443 6052 6452
rect 6000 6409 6009 6443
rect 6009 6409 6043 6443
rect 6043 6409 6052 6443
rect 6000 6400 6052 6409
rect 7656 6400 7708 6452
rect 6644 6332 6696 6384
rect 4344 6239 4396 6248
rect 4344 6205 4353 6239
rect 4353 6205 4387 6239
rect 4387 6205 4396 6239
rect 4344 6196 4396 6205
rect 7564 6264 7616 6316
rect 7656 6307 7708 6316
rect 7656 6273 7665 6307
rect 7665 6273 7699 6307
rect 7699 6273 7708 6307
rect 7656 6264 7708 6273
rect 8208 6400 8260 6452
rect 8668 6443 8720 6452
rect 8668 6409 8677 6443
rect 8677 6409 8711 6443
rect 8711 6409 8720 6443
rect 8668 6400 8720 6409
rect 8392 6307 8444 6316
rect 8392 6273 8406 6307
rect 8406 6273 8440 6307
rect 8440 6273 8444 6307
rect 8392 6264 8444 6273
rect 2780 6060 2832 6112
rect 3424 6103 3476 6112
rect 3424 6069 3433 6103
rect 3433 6069 3467 6103
rect 3467 6069 3476 6103
rect 3424 6060 3476 6069
rect 4528 6060 4580 6112
rect 5080 6103 5132 6112
rect 5080 6069 5089 6103
rect 5089 6069 5123 6103
rect 5123 6069 5132 6103
rect 5080 6060 5132 6069
rect 7932 6128 7984 6180
rect 8484 6128 8536 6180
rect 6828 6060 6880 6112
rect 7472 6060 7524 6112
rect 7564 6103 7616 6112
rect 7564 6069 7573 6103
rect 7573 6069 7607 6103
rect 7607 6069 7616 6103
rect 7564 6060 7616 6069
rect 7656 6060 7708 6112
rect 1985 5958 2037 6010
rect 2049 5958 2101 6010
rect 2113 5958 2165 6010
rect 2177 5958 2229 6010
rect 2241 5958 2293 6010
rect 4055 5958 4107 6010
rect 4119 5958 4171 6010
rect 4183 5958 4235 6010
rect 4247 5958 4299 6010
rect 4311 5958 4363 6010
rect 6125 5958 6177 6010
rect 6189 5958 6241 6010
rect 6253 5958 6305 6010
rect 6317 5958 6369 6010
rect 6381 5958 6433 6010
rect 8195 5958 8247 6010
rect 8259 5958 8311 6010
rect 8323 5958 8375 6010
rect 8387 5958 8439 6010
rect 8451 5958 8503 6010
rect 1860 5856 1912 5908
rect 2780 5899 2832 5908
rect 2780 5865 2789 5899
rect 2789 5865 2823 5899
rect 2823 5865 2832 5899
rect 2780 5856 2832 5865
rect 3424 5856 3476 5908
rect 5356 5856 5408 5908
rect 6644 5856 6696 5908
rect 7196 5856 7248 5908
rect 2136 5720 2188 5772
rect 2320 5720 2372 5772
rect 7932 5856 7984 5908
rect 8668 5899 8720 5908
rect 8668 5865 8677 5899
rect 8677 5865 8711 5899
rect 8711 5865 8720 5899
rect 8668 5856 8720 5865
rect 1584 5652 1636 5704
rect 1768 5695 1820 5704
rect 1768 5661 1777 5695
rect 1777 5661 1811 5695
rect 1811 5661 1820 5695
rect 1768 5652 1820 5661
rect 2228 5652 2280 5704
rect 3148 5652 3200 5704
rect 3884 5652 3936 5704
rect 4068 5695 4120 5704
rect 4068 5661 4077 5695
rect 4077 5661 4111 5695
rect 4111 5661 4120 5695
rect 4068 5652 4120 5661
rect 1952 5516 2004 5568
rect 4436 5652 4488 5704
rect 5080 5695 5132 5704
rect 5080 5661 5089 5695
rect 5089 5661 5123 5695
rect 5123 5661 5132 5695
rect 5080 5652 5132 5661
rect 5816 5584 5868 5636
rect 7656 5695 7708 5704
rect 7656 5661 7665 5695
rect 7665 5661 7699 5695
rect 7699 5661 7708 5695
rect 7656 5652 7708 5661
rect 7564 5584 7616 5636
rect 8024 5652 8076 5704
rect 4528 5516 4580 5568
rect 8116 5516 8168 5568
rect 2645 5414 2697 5466
rect 2709 5414 2761 5466
rect 2773 5414 2825 5466
rect 2837 5414 2889 5466
rect 2901 5414 2953 5466
rect 4715 5414 4767 5466
rect 4779 5414 4831 5466
rect 4843 5414 4895 5466
rect 4907 5414 4959 5466
rect 4971 5414 5023 5466
rect 6785 5414 6837 5466
rect 6849 5414 6901 5466
rect 6913 5414 6965 5466
rect 6977 5414 7029 5466
rect 7041 5414 7093 5466
rect 8855 5414 8907 5466
rect 8919 5414 8971 5466
rect 8983 5414 9035 5466
rect 9047 5414 9099 5466
rect 9111 5414 9163 5466
rect 1400 5312 1452 5364
rect 1768 5355 1820 5364
rect 1768 5321 1777 5355
rect 1777 5321 1811 5355
rect 1811 5321 1820 5355
rect 1768 5312 1820 5321
rect 2320 5312 2372 5364
rect 5080 5312 5132 5364
rect 8024 5355 8076 5364
rect 8024 5321 8033 5355
rect 8033 5321 8067 5355
rect 8067 5321 8076 5355
rect 8024 5312 8076 5321
rect 1584 5176 1636 5228
rect 1952 5219 2004 5228
rect 1952 5185 1961 5219
rect 1961 5185 1995 5219
rect 1995 5185 2004 5219
rect 1952 5176 2004 5185
rect 2872 5219 2924 5228
rect 2872 5185 2881 5219
rect 2881 5185 2915 5219
rect 2915 5185 2924 5219
rect 2872 5176 2924 5185
rect 4436 5176 4488 5228
rect 2136 5108 2188 5160
rect 4528 5151 4580 5160
rect 4528 5117 4537 5151
rect 4537 5117 4571 5151
rect 4571 5117 4580 5151
rect 4528 5108 4580 5117
rect 5356 5219 5408 5228
rect 5356 5185 5365 5219
rect 5365 5185 5399 5219
rect 5399 5185 5408 5219
rect 5356 5176 5408 5185
rect 5632 5176 5684 5228
rect 8208 5176 8260 5228
rect 3424 5040 3476 5092
rect 4068 5040 4120 5092
rect 5172 5040 5224 5092
rect 7564 5151 7616 5160
rect 7564 5117 7573 5151
rect 7573 5117 7607 5151
rect 7607 5117 7616 5151
rect 7564 5108 7616 5117
rect 7748 5151 7800 5160
rect 7748 5117 7757 5151
rect 7757 5117 7791 5151
rect 7791 5117 7800 5151
rect 7748 5108 7800 5117
rect 7840 5151 7892 5160
rect 7840 5117 7849 5151
rect 7849 5117 7883 5151
rect 7883 5117 7892 5151
rect 7840 5108 7892 5117
rect 8024 5108 8076 5160
rect 9036 5151 9088 5160
rect 9036 5117 9045 5151
rect 9045 5117 9079 5151
rect 9079 5117 9088 5151
rect 9036 5108 9088 5117
rect 3056 5015 3108 5024
rect 3056 4981 3065 5015
rect 3065 4981 3099 5015
rect 3099 4981 3108 5015
rect 3056 4972 3108 4981
rect 4896 5015 4948 5024
rect 4896 4981 4905 5015
rect 4905 4981 4939 5015
rect 4939 4981 4948 5015
rect 4896 4972 4948 4981
rect 5448 4972 5500 5024
rect 6552 4972 6604 5024
rect 7196 4972 7248 5024
rect 1985 4870 2037 4922
rect 2049 4870 2101 4922
rect 2113 4870 2165 4922
rect 2177 4870 2229 4922
rect 2241 4870 2293 4922
rect 4055 4870 4107 4922
rect 4119 4870 4171 4922
rect 4183 4870 4235 4922
rect 4247 4870 4299 4922
rect 4311 4870 4363 4922
rect 6125 4870 6177 4922
rect 6189 4870 6241 4922
rect 6253 4870 6305 4922
rect 6317 4870 6369 4922
rect 6381 4870 6433 4922
rect 8195 4870 8247 4922
rect 8259 4870 8311 4922
rect 8323 4870 8375 4922
rect 8387 4870 8439 4922
rect 8451 4870 8503 4922
rect 2872 4768 2924 4820
rect 4896 4768 4948 4820
rect 5448 4811 5500 4820
rect 5448 4777 5457 4811
rect 5457 4777 5491 4811
rect 5491 4777 5500 4811
rect 5448 4768 5500 4777
rect 2964 4700 3016 4752
rect 2596 4632 2648 4684
rect 5540 4700 5592 4752
rect 7104 4768 7156 4820
rect 7196 4811 7248 4820
rect 7196 4777 7205 4811
rect 7205 4777 7239 4811
rect 7239 4777 7248 4811
rect 7196 4768 7248 4777
rect 7840 4768 7892 4820
rect 940 4564 992 4616
rect 1584 4564 1636 4616
rect 3056 4564 3108 4616
rect 3884 4564 3936 4616
rect 4068 4607 4120 4616
rect 4068 4573 4077 4607
rect 4077 4573 4111 4607
rect 4111 4573 4120 4607
rect 4068 4564 4120 4573
rect 5080 4564 5132 4616
rect 3792 4471 3844 4480
rect 3792 4437 3801 4471
rect 3801 4437 3835 4471
rect 3835 4437 3844 4471
rect 3792 4428 3844 4437
rect 5356 4496 5408 4548
rect 7656 4700 7708 4752
rect 7288 4675 7340 4684
rect 7288 4641 7297 4675
rect 7297 4641 7331 4675
rect 7331 4641 7340 4675
rect 7288 4632 7340 4641
rect 6644 4564 6696 4616
rect 8024 4700 8076 4752
rect 8116 4607 8168 4616
rect 8116 4573 8125 4607
rect 8125 4573 8159 4607
rect 8159 4573 8168 4607
rect 8116 4564 8168 4573
rect 5172 4471 5224 4480
rect 5172 4437 5181 4471
rect 5181 4437 5215 4471
rect 5215 4437 5224 4471
rect 5172 4428 5224 4437
rect 5632 4428 5684 4480
rect 5724 4428 5776 4480
rect 7196 4428 7248 4480
rect 2645 4326 2697 4378
rect 2709 4326 2761 4378
rect 2773 4326 2825 4378
rect 2837 4326 2889 4378
rect 2901 4326 2953 4378
rect 4715 4326 4767 4378
rect 4779 4326 4831 4378
rect 4843 4326 4895 4378
rect 4907 4326 4959 4378
rect 4971 4326 5023 4378
rect 6785 4326 6837 4378
rect 6849 4326 6901 4378
rect 6913 4326 6965 4378
rect 6977 4326 7029 4378
rect 7041 4326 7093 4378
rect 8855 4326 8907 4378
rect 8919 4326 8971 4378
rect 8983 4326 9035 4378
rect 9047 4326 9099 4378
rect 9111 4326 9163 4378
rect 1676 4131 1728 4140
rect 1676 4097 1685 4131
rect 1685 4097 1719 4131
rect 1719 4097 1728 4131
rect 1676 4088 1728 4097
rect 1860 4131 1912 4140
rect 1860 4097 1869 4131
rect 1869 4097 1903 4131
rect 1903 4097 1912 4131
rect 1860 4088 1912 4097
rect 3424 4088 3476 4140
rect 7288 4224 7340 4276
rect 3792 4088 3844 4140
rect 4436 4088 4488 4140
rect 6552 4088 6604 4140
rect 3976 4020 4028 4072
rect 7288 4063 7340 4072
rect 7288 4029 7297 4063
rect 7297 4029 7331 4063
rect 7331 4029 7340 4063
rect 7288 4020 7340 4029
rect 7748 4020 7800 4072
rect 3424 3884 3476 3936
rect 7380 3884 7432 3936
rect 7748 3884 7800 3936
rect 1985 3782 2037 3834
rect 2049 3782 2101 3834
rect 2113 3782 2165 3834
rect 2177 3782 2229 3834
rect 2241 3782 2293 3834
rect 4055 3782 4107 3834
rect 4119 3782 4171 3834
rect 4183 3782 4235 3834
rect 4247 3782 4299 3834
rect 4311 3782 4363 3834
rect 6125 3782 6177 3834
rect 6189 3782 6241 3834
rect 6253 3782 6305 3834
rect 6317 3782 6369 3834
rect 6381 3782 6433 3834
rect 8195 3782 8247 3834
rect 8259 3782 8311 3834
rect 8323 3782 8375 3834
rect 8387 3782 8439 3834
rect 8451 3782 8503 3834
rect 1584 3723 1636 3732
rect 1584 3689 1593 3723
rect 1593 3689 1627 3723
rect 1627 3689 1636 3723
rect 1584 3680 1636 3689
rect 1860 3680 1912 3732
rect 3976 3680 4028 3732
rect 5080 3723 5132 3732
rect 5080 3689 5089 3723
rect 5089 3689 5123 3723
rect 5123 3689 5132 3723
rect 5080 3680 5132 3689
rect 5540 3680 5592 3732
rect 2136 3587 2188 3596
rect 2136 3553 2145 3587
rect 2145 3553 2179 3587
rect 2179 3553 2188 3587
rect 2136 3544 2188 3553
rect 4344 3655 4396 3664
rect 4344 3621 4353 3655
rect 4353 3621 4387 3655
rect 4387 3621 4396 3655
rect 4344 3612 4396 3621
rect 2412 3544 2464 3596
rect 940 3408 992 3460
rect 2228 3519 2280 3528
rect 2228 3485 2237 3519
rect 2237 3485 2271 3519
rect 2271 3485 2280 3519
rect 2228 3476 2280 3485
rect 3240 3476 3292 3528
rect 4436 3476 4488 3528
rect 4620 3519 4672 3528
rect 4620 3485 4629 3519
rect 4629 3485 4663 3519
rect 4663 3485 4672 3519
rect 4620 3476 4672 3485
rect 7380 3587 7432 3596
rect 7380 3553 7389 3587
rect 7389 3553 7423 3587
rect 7423 3553 7432 3587
rect 7380 3544 7432 3553
rect 7472 3544 7524 3596
rect 3148 3451 3200 3460
rect 3148 3417 3157 3451
rect 3157 3417 3191 3451
rect 3191 3417 3200 3451
rect 3148 3408 3200 3417
rect 3332 3451 3384 3460
rect 3332 3417 3341 3451
rect 3341 3417 3375 3451
rect 3375 3417 3384 3451
rect 3332 3408 3384 3417
rect 5356 3519 5408 3528
rect 5356 3485 5365 3519
rect 5365 3485 5399 3519
rect 5399 3485 5408 3519
rect 5356 3476 5408 3485
rect 5540 3519 5592 3528
rect 5540 3485 5549 3519
rect 5549 3485 5583 3519
rect 5583 3485 5592 3519
rect 5540 3476 5592 3485
rect 7196 3476 7248 3528
rect 8668 3519 8720 3528
rect 8668 3485 8677 3519
rect 8677 3485 8711 3519
rect 8711 3485 8720 3519
rect 8668 3476 8720 3485
rect 3056 3340 3108 3392
rect 5080 3340 5132 3392
rect 7748 3340 7800 3392
rect 2645 3238 2697 3290
rect 2709 3238 2761 3290
rect 2773 3238 2825 3290
rect 2837 3238 2889 3290
rect 2901 3238 2953 3290
rect 4715 3238 4767 3290
rect 4779 3238 4831 3290
rect 4843 3238 4895 3290
rect 4907 3238 4959 3290
rect 4971 3238 5023 3290
rect 6785 3238 6837 3290
rect 6849 3238 6901 3290
rect 6913 3238 6965 3290
rect 6977 3238 7029 3290
rect 7041 3238 7093 3290
rect 8855 3238 8907 3290
rect 8919 3238 8971 3290
rect 8983 3238 9035 3290
rect 9047 3238 9099 3290
rect 9111 3238 9163 3290
rect 1492 3136 1544 3188
rect 1400 3068 1452 3120
rect 2228 3136 2280 3188
rect 3148 3136 3200 3188
rect 3332 3136 3384 3188
rect 3424 3179 3476 3188
rect 3424 3145 3433 3179
rect 3433 3145 3467 3179
rect 3467 3145 3476 3179
rect 3424 3136 3476 3145
rect 4344 3136 4396 3188
rect 4436 3136 4488 3188
rect 1860 3043 1912 3052
rect 1860 3009 1869 3043
rect 1869 3009 1903 3043
rect 1903 3009 1912 3043
rect 1860 3000 1912 3009
rect 2136 3068 2188 3120
rect 3056 3068 3108 3120
rect 2320 3043 2372 3052
rect 2320 3009 2329 3043
rect 2329 3009 2363 3043
rect 2363 3009 2372 3043
rect 2320 3000 2372 3009
rect 1860 2864 1912 2916
rect 3056 2932 3108 2984
rect 4620 3000 4672 3052
rect 5540 3136 5592 3188
rect 7288 3136 7340 3188
rect 7380 3136 7432 3188
rect 7564 3136 7616 3188
rect 8576 3136 8628 3188
rect 5080 3043 5132 3052
rect 5080 3009 5089 3043
rect 5089 3009 5123 3043
rect 5123 3009 5132 3043
rect 5080 3000 5132 3009
rect 5448 3000 5500 3052
rect 5632 3043 5684 3052
rect 5632 3009 5641 3043
rect 5641 3009 5675 3043
rect 5675 3009 5684 3043
rect 5632 3000 5684 3009
rect 6460 3000 6512 3052
rect 7196 3000 7248 3052
rect 4436 2932 4488 2984
rect 2136 2796 2188 2848
rect 5356 2864 5408 2916
rect 5724 2796 5776 2848
rect 7564 3043 7616 3052
rect 7564 3009 7573 3043
rect 7573 3009 7607 3043
rect 7607 3009 7616 3043
rect 7564 3000 7616 3009
rect 7932 3043 7984 3052
rect 7932 3009 7941 3043
rect 7941 3009 7975 3043
rect 7975 3009 7984 3043
rect 7932 3000 7984 3009
rect 8116 3000 8168 3052
rect 9404 3000 9456 3052
rect 6736 2796 6788 2848
rect 7380 2839 7432 2848
rect 7380 2805 7389 2839
rect 7389 2805 7423 2839
rect 7423 2805 7432 2839
rect 7380 2796 7432 2805
rect 1985 2694 2037 2746
rect 2049 2694 2101 2746
rect 2113 2694 2165 2746
rect 2177 2694 2229 2746
rect 2241 2694 2293 2746
rect 4055 2694 4107 2746
rect 4119 2694 4171 2746
rect 4183 2694 4235 2746
rect 4247 2694 4299 2746
rect 4311 2694 4363 2746
rect 6125 2694 6177 2746
rect 6189 2694 6241 2746
rect 6253 2694 6305 2746
rect 6317 2694 6369 2746
rect 6381 2694 6433 2746
rect 8195 2694 8247 2746
rect 8259 2694 8311 2746
rect 8323 2694 8375 2746
rect 8387 2694 8439 2746
rect 8451 2694 8503 2746
rect 3516 2592 3568 2644
rect 4436 2592 4488 2644
rect 5632 2592 5684 2644
rect 6000 2635 6052 2644
rect 6000 2601 6009 2635
rect 6009 2601 6043 2635
rect 6043 2601 6052 2635
rect 6000 2592 6052 2601
rect 6644 2592 6696 2644
rect 7564 2592 7616 2644
rect 6736 2524 6788 2576
rect 1308 2456 1360 2508
rect 1216 2388 1268 2440
rect 5448 2431 5500 2440
rect 5448 2397 5457 2431
rect 5457 2397 5491 2431
rect 5491 2397 5500 2431
rect 5448 2388 5500 2397
rect 5540 2431 5592 2440
rect 5540 2397 5549 2431
rect 5549 2397 5583 2431
rect 5583 2397 5592 2431
rect 5540 2388 5592 2397
rect 5816 2388 5868 2440
rect 20 2320 72 2372
rect 3240 2320 3292 2372
rect 5724 2363 5776 2372
rect 5724 2329 5733 2363
rect 5733 2329 5767 2363
rect 5767 2329 5776 2363
rect 5724 2320 5776 2329
rect 7196 2456 7248 2508
rect 7564 2431 7616 2440
rect 7564 2397 7573 2431
rect 7573 2397 7607 2431
rect 7607 2397 7616 2431
rect 7564 2388 7616 2397
rect 5632 2252 5684 2304
rect 7380 2320 7432 2372
rect 6552 2252 6604 2304
rect 7748 2320 7800 2372
rect 7932 2320 7984 2372
rect 10324 2320 10376 2372
rect 2645 2150 2697 2202
rect 2709 2150 2761 2202
rect 2773 2150 2825 2202
rect 2837 2150 2889 2202
rect 2901 2150 2953 2202
rect 4715 2150 4767 2202
rect 4779 2150 4831 2202
rect 4843 2150 4895 2202
rect 4907 2150 4959 2202
rect 4971 2150 5023 2202
rect 6785 2150 6837 2202
rect 6849 2150 6901 2202
rect 6913 2150 6965 2202
rect 6977 2150 7029 2202
rect 7041 2150 7093 2202
rect 8855 2150 8907 2202
rect 8919 2150 8971 2202
rect 8983 2150 9035 2202
rect 9047 2150 9099 2202
rect 9111 2150 9163 2202
rect 5724 2048 5776 2100
rect 7748 2048 7800 2100
<< metal2 >>
rect 1306 11911 1362 12711
rect 2594 11911 2650 12711
rect 4526 12050 4582 12711
rect 6458 12050 6514 12711
rect 4526 12022 4660 12050
rect 2778 11928 2834 11937
rect 1320 10062 1348 11911
rect 1985 10364 2293 10373
rect 1985 10362 1991 10364
rect 2047 10362 2071 10364
rect 2127 10362 2151 10364
rect 2207 10362 2231 10364
rect 2287 10362 2293 10364
rect 2047 10310 2049 10362
rect 2229 10310 2231 10362
rect 1985 10308 1991 10310
rect 2047 10308 2071 10310
rect 2127 10308 2151 10310
rect 2207 10308 2231 10310
rect 2287 10308 2293 10310
rect 1985 10299 2293 10308
rect 1398 10160 1454 10169
rect 1398 10095 1454 10104
rect 1308 10056 1360 10062
rect 1308 9998 1360 10004
rect 1412 9586 1440 10095
rect 2608 10062 2636 11911
rect 4526 11911 4582 12022
rect 2778 11863 2834 11872
rect 2792 10198 2820 11863
rect 4055 10364 4363 10373
rect 4055 10362 4061 10364
rect 4117 10362 4141 10364
rect 4197 10362 4221 10364
rect 4277 10362 4301 10364
rect 4357 10362 4363 10364
rect 4117 10310 4119 10362
rect 4299 10310 4301 10362
rect 4055 10308 4061 10310
rect 4117 10308 4141 10310
rect 4197 10308 4221 10310
rect 4277 10308 4301 10310
rect 4357 10308 4363 10310
rect 4055 10299 4363 10308
rect 4632 10266 4660 12022
rect 6458 12022 6776 12050
rect 6458 11911 6514 12022
rect 6125 10364 6433 10373
rect 6125 10362 6131 10364
rect 6187 10362 6211 10364
rect 6267 10362 6291 10364
rect 6347 10362 6371 10364
rect 6427 10362 6433 10364
rect 6187 10310 6189 10362
rect 6369 10310 6371 10362
rect 6125 10308 6131 10310
rect 6187 10308 6211 10310
rect 6267 10308 6291 10310
rect 6347 10308 6371 10310
rect 6427 10308 6433 10310
rect 6125 10299 6433 10308
rect 6748 10266 6776 12022
rect 7746 11911 7802 12711
rect 9678 11911 9734 12711
rect 4620 10260 4672 10266
rect 4620 10202 4672 10208
rect 6736 10260 6788 10266
rect 6736 10202 6788 10208
rect 2780 10192 2832 10198
rect 2780 10134 2832 10140
rect 7760 10062 7788 11911
rect 9310 11656 9366 11665
rect 9310 11591 9366 11600
rect 8195 10364 8503 10373
rect 8195 10362 8201 10364
rect 8257 10362 8281 10364
rect 8337 10362 8361 10364
rect 8417 10362 8441 10364
rect 8497 10362 8503 10364
rect 8257 10310 8259 10362
rect 8439 10310 8441 10362
rect 8195 10308 8201 10310
rect 8257 10308 8281 10310
rect 8337 10308 8361 10310
rect 8417 10308 8441 10310
rect 8497 10308 8503 10310
rect 8195 10299 8503 10308
rect 2596 10056 2648 10062
rect 2596 9998 2648 10004
rect 4160 10056 4212 10062
rect 4160 9998 4212 10004
rect 7748 10056 7800 10062
rect 7748 9998 7800 10004
rect 8484 10056 8536 10062
rect 8668 10056 8720 10062
rect 8536 10016 8616 10044
rect 8484 9998 8536 10004
rect 1676 9988 1728 9994
rect 2504 9988 2556 9994
rect 1728 9948 1900 9976
rect 1676 9930 1728 9936
rect 1400 9580 1452 9586
rect 1400 9522 1452 9528
rect 1676 9512 1728 9518
rect 1676 9454 1728 9460
rect 1400 9376 1452 9382
rect 1400 9318 1452 9324
rect 940 8968 992 8974
rect 938 8936 940 8945
rect 992 8936 994 8945
rect 938 8871 994 8880
rect 1412 5370 1440 9318
rect 1688 7528 1716 9454
rect 1768 9444 1820 9450
rect 1768 9386 1820 9392
rect 1780 8974 1808 9386
rect 1768 8968 1820 8974
rect 1768 8910 1820 8916
rect 1768 8424 1820 8430
rect 1768 8366 1820 8372
rect 1780 8090 1808 8366
rect 1768 8084 1820 8090
rect 1768 8026 1820 8032
rect 1596 7500 1716 7528
rect 1492 7200 1544 7206
rect 1492 7142 1544 7148
rect 1504 6905 1532 7142
rect 1490 6896 1546 6905
rect 1490 6831 1546 6840
rect 1596 5794 1624 7500
rect 1768 7404 1820 7410
rect 1768 7346 1820 7352
rect 1780 7154 1808 7346
rect 1504 5766 1624 5794
rect 1688 7126 1808 7154
rect 1400 5364 1452 5370
rect 1400 5306 1452 5312
rect 938 4856 994 4865
rect 938 4791 994 4800
rect 952 4622 980 4791
rect 940 4616 992 4622
rect 940 4558 992 4564
rect 938 3496 994 3505
rect 938 3431 940 3440
rect 992 3431 994 3440
rect 940 3402 992 3408
rect 1412 3126 1440 5306
rect 1504 3194 1532 5766
rect 1584 5704 1636 5710
rect 1584 5646 1636 5652
rect 1596 5234 1624 5646
rect 1584 5228 1636 5234
rect 1584 5170 1636 5176
rect 1596 4622 1624 5170
rect 1584 4616 1636 4622
rect 1584 4558 1636 4564
rect 1596 3738 1624 4558
rect 1688 4146 1716 7126
rect 1872 6798 1900 9948
rect 2504 9930 2556 9936
rect 2320 9580 2372 9586
rect 2320 9522 2372 9528
rect 2332 9466 2360 9522
rect 2332 9438 2452 9466
rect 1985 9276 2293 9285
rect 1985 9274 1991 9276
rect 2047 9274 2071 9276
rect 2127 9274 2151 9276
rect 2207 9274 2231 9276
rect 2287 9274 2293 9276
rect 2047 9222 2049 9274
rect 2229 9222 2231 9274
rect 1985 9220 1991 9222
rect 2047 9220 2071 9222
rect 2127 9220 2151 9222
rect 2207 9220 2231 9222
rect 2287 9220 2293 9222
rect 1985 9211 2293 9220
rect 2424 8974 2452 9438
rect 2412 8968 2464 8974
rect 2412 8910 2464 8916
rect 2424 8566 2452 8910
rect 2412 8560 2464 8566
rect 2412 8502 2464 8508
rect 2412 8288 2464 8294
rect 2412 8230 2464 8236
rect 1985 8188 2293 8197
rect 1985 8186 1991 8188
rect 2047 8186 2071 8188
rect 2127 8186 2151 8188
rect 2207 8186 2231 8188
rect 2287 8186 2293 8188
rect 2047 8134 2049 8186
rect 2229 8134 2231 8186
rect 1985 8132 1991 8134
rect 2047 8132 2071 8134
rect 2127 8132 2151 8134
rect 2207 8132 2231 8134
rect 2287 8132 2293 8134
rect 1985 8123 2293 8132
rect 2424 7886 2452 8230
rect 2412 7880 2464 7886
rect 2412 7822 2464 7828
rect 2320 7812 2372 7818
rect 2320 7754 2372 7760
rect 2332 7546 2360 7754
rect 2320 7540 2372 7546
rect 2320 7482 2372 7488
rect 2424 7410 2452 7822
rect 2412 7404 2464 7410
rect 2412 7346 2464 7352
rect 2412 7200 2464 7206
rect 2412 7142 2464 7148
rect 1985 7100 2293 7109
rect 1985 7098 1991 7100
rect 2047 7098 2071 7100
rect 2127 7098 2151 7100
rect 2207 7098 2231 7100
rect 2287 7098 2293 7100
rect 2047 7046 2049 7098
rect 2229 7046 2231 7098
rect 1985 7044 1991 7046
rect 2047 7044 2071 7046
rect 2127 7044 2151 7046
rect 2207 7044 2231 7046
rect 2287 7044 2293 7046
rect 1985 7035 2293 7044
rect 2136 6996 2188 7002
rect 2136 6938 2188 6944
rect 1860 6792 1912 6798
rect 1860 6734 1912 6740
rect 1872 6458 1900 6734
rect 1860 6452 1912 6458
rect 1860 6394 1912 6400
rect 1872 5914 1900 6394
rect 2148 6390 2176 6938
rect 2424 6866 2452 7142
rect 2320 6860 2372 6866
rect 2320 6802 2372 6808
rect 2412 6860 2464 6866
rect 2412 6802 2464 6808
rect 2136 6384 2188 6390
rect 2136 6326 2188 6332
rect 1985 6012 2293 6021
rect 1985 6010 1991 6012
rect 2047 6010 2071 6012
rect 2127 6010 2151 6012
rect 2207 6010 2231 6012
rect 2287 6010 2293 6012
rect 2047 5958 2049 6010
rect 2229 5958 2231 6010
rect 1985 5956 1991 5958
rect 2047 5956 2071 5958
rect 2127 5956 2151 5958
rect 2207 5956 2231 5958
rect 2287 5956 2293 5958
rect 1985 5947 2293 5956
rect 1860 5908 1912 5914
rect 1860 5850 1912 5856
rect 2332 5778 2360 6802
rect 2424 6322 2452 6802
rect 2412 6316 2464 6322
rect 2412 6258 2464 6264
rect 2136 5772 2188 5778
rect 2136 5714 2188 5720
rect 2320 5772 2372 5778
rect 2320 5714 2372 5720
rect 1768 5704 1820 5710
rect 1768 5646 1820 5652
rect 1780 5370 1808 5646
rect 1952 5568 2004 5574
rect 1952 5510 2004 5516
rect 1768 5364 1820 5370
rect 1768 5306 1820 5312
rect 1964 5234 1992 5510
rect 1952 5228 2004 5234
rect 1952 5170 2004 5176
rect 1964 5012 1992 5170
rect 2148 5166 2176 5714
rect 2228 5704 2280 5710
rect 2228 5646 2280 5652
rect 2240 5250 2268 5646
rect 2332 5370 2360 5714
rect 2320 5364 2372 5370
rect 2320 5306 2372 5312
rect 2240 5222 2452 5250
rect 2136 5160 2188 5166
rect 2136 5102 2188 5108
rect 1964 4984 2360 5012
rect 1985 4924 2293 4933
rect 1985 4922 1991 4924
rect 2047 4922 2071 4924
rect 2127 4922 2151 4924
rect 2207 4922 2231 4924
rect 2287 4922 2293 4924
rect 2047 4870 2049 4922
rect 2229 4870 2231 4922
rect 1985 4868 1991 4870
rect 2047 4868 2071 4870
rect 2127 4868 2151 4870
rect 2207 4868 2231 4870
rect 2287 4868 2293 4870
rect 1985 4859 2293 4868
rect 1676 4140 1728 4146
rect 1676 4082 1728 4088
rect 1860 4140 1912 4146
rect 1860 4082 1912 4088
rect 1872 3738 1900 4082
rect 1985 3836 2293 3845
rect 1985 3834 1991 3836
rect 2047 3834 2071 3836
rect 2127 3834 2151 3836
rect 2207 3834 2231 3836
rect 2287 3834 2293 3836
rect 2047 3782 2049 3834
rect 2229 3782 2231 3834
rect 1985 3780 1991 3782
rect 2047 3780 2071 3782
rect 2127 3780 2151 3782
rect 2207 3780 2231 3782
rect 2287 3780 2293 3782
rect 1985 3771 2293 3780
rect 1584 3732 1636 3738
rect 1584 3674 1636 3680
rect 1860 3732 1912 3738
rect 1860 3674 1912 3680
rect 2136 3596 2188 3602
rect 2136 3538 2188 3544
rect 1492 3188 1544 3194
rect 1492 3130 1544 3136
rect 2148 3126 2176 3538
rect 2228 3528 2280 3534
rect 2228 3470 2280 3476
rect 2240 3194 2268 3470
rect 2228 3188 2280 3194
rect 2228 3130 2280 3136
rect 1400 3120 1452 3126
rect 1400 3062 1452 3068
rect 2136 3120 2188 3126
rect 2136 3062 2188 3068
rect 1860 3052 1912 3058
rect 1860 2994 1912 3000
rect 1872 2922 1900 2994
rect 1860 2916 1912 2922
rect 1860 2858 1912 2864
rect 2148 2854 2176 3062
rect 2332 3058 2360 4984
rect 2424 3602 2452 5222
rect 2516 4672 2544 9930
rect 2645 9820 2953 9829
rect 2645 9818 2651 9820
rect 2707 9818 2731 9820
rect 2787 9818 2811 9820
rect 2867 9818 2891 9820
rect 2947 9818 2953 9820
rect 2707 9766 2709 9818
rect 2889 9766 2891 9818
rect 2645 9764 2651 9766
rect 2707 9764 2731 9766
rect 2787 9764 2811 9766
rect 2867 9764 2891 9766
rect 2947 9764 2953 9766
rect 2645 9755 2953 9764
rect 3238 9616 3294 9625
rect 2688 9580 2740 9586
rect 2688 9522 2740 9528
rect 3056 9580 3108 9586
rect 3238 9551 3240 9560
rect 3056 9522 3108 9528
rect 3292 9551 3294 9560
rect 4068 9580 4120 9586
rect 3240 9522 3292 9528
rect 4068 9522 4120 9528
rect 2596 9376 2648 9382
rect 2596 9318 2648 9324
rect 2608 9178 2636 9318
rect 2700 9178 2728 9522
rect 2596 9172 2648 9178
rect 2596 9114 2648 9120
rect 2688 9172 2740 9178
rect 2688 9114 2740 9120
rect 2645 8732 2953 8741
rect 2645 8730 2651 8732
rect 2707 8730 2731 8732
rect 2787 8730 2811 8732
rect 2867 8730 2891 8732
rect 2947 8730 2953 8732
rect 2707 8678 2709 8730
rect 2889 8678 2891 8730
rect 2645 8676 2651 8678
rect 2707 8676 2731 8678
rect 2787 8676 2811 8678
rect 2867 8676 2891 8678
rect 2947 8676 2953 8678
rect 2645 8667 2953 8676
rect 3068 8566 3096 9522
rect 3792 9512 3844 9518
rect 3792 9454 3844 9460
rect 3976 9512 4028 9518
rect 3976 9454 4028 9460
rect 3240 9376 3292 9382
rect 3240 9318 3292 9324
rect 3252 9178 3280 9318
rect 3240 9172 3292 9178
rect 3240 9114 3292 9120
rect 3148 9104 3200 9110
rect 3148 9046 3200 9052
rect 3056 8560 3108 8566
rect 3056 8502 3108 8508
rect 2780 8288 2832 8294
rect 2780 8230 2832 8236
rect 2792 7954 2820 8230
rect 2780 7948 2832 7954
rect 2780 7890 2832 7896
rect 2645 7644 2953 7653
rect 2645 7642 2651 7644
rect 2707 7642 2731 7644
rect 2787 7642 2811 7644
rect 2867 7642 2891 7644
rect 2947 7642 2953 7644
rect 2707 7590 2709 7642
rect 2889 7590 2891 7642
rect 2645 7588 2651 7590
rect 2707 7588 2731 7590
rect 2787 7588 2811 7590
rect 2867 7588 2891 7590
rect 2947 7588 2953 7590
rect 2645 7579 2953 7588
rect 2688 7404 2740 7410
rect 2688 7346 2740 7352
rect 2700 7002 2728 7346
rect 3068 7206 3096 8502
rect 3056 7200 3108 7206
rect 3056 7142 3108 7148
rect 2688 6996 2740 7002
rect 2688 6938 2740 6944
rect 2645 6556 2953 6565
rect 2645 6554 2651 6556
rect 2707 6554 2731 6556
rect 2787 6554 2811 6556
rect 2867 6554 2891 6556
rect 2947 6554 2953 6556
rect 2707 6502 2709 6554
rect 2889 6502 2891 6554
rect 2645 6500 2651 6502
rect 2707 6500 2731 6502
rect 2787 6500 2811 6502
rect 2867 6500 2891 6502
rect 2947 6500 2953 6502
rect 2645 6491 2953 6500
rect 2780 6112 2832 6118
rect 2780 6054 2832 6060
rect 2792 5914 2820 6054
rect 2780 5908 2832 5914
rect 2780 5850 2832 5856
rect 2645 5468 2953 5477
rect 2645 5466 2651 5468
rect 2707 5466 2731 5468
rect 2787 5466 2811 5468
rect 2867 5466 2891 5468
rect 2947 5466 2953 5468
rect 2707 5414 2709 5466
rect 2889 5414 2891 5466
rect 2645 5412 2651 5414
rect 2707 5412 2731 5414
rect 2787 5412 2811 5414
rect 2867 5412 2891 5414
rect 2947 5412 2953 5414
rect 2645 5403 2953 5412
rect 3068 5386 3096 7142
rect 3160 5710 3188 9046
rect 3804 8922 3832 9454
rect 3988 9110 4016 9454
rect 4080 9382 4108 9522
rect 4172 9450 4200 9998
rect 5080 9988 5132 9994
rect 5080 9930 5132 9936
rect 7288 9988 7340 9994
rect 7288 9930 7340 9936
rect 4715 9820 5023 9829
rect 4715 9818 4721 9820
rect 4777 9818 4801 9820
rect 4857 9818 4881 9820
rect 4937 9818 4961 9820
rect 5017 9818 5023 9820
rect 4777 9766 4779 9818
rect 4959 9766 4961 9818
rect 4715 9764 4721 9766
rect 4777 9764 4801 9766
rect 4857 9764 4881 9766
rect 4937 9764 4961 9766
rect 5017 9764 5023 9766
rect 4715 9755 5023 9764
rect 5092 9722 5120 9930
rect 6644 9920 6696 9926
rect 6644 9862 6696 9868
rect 5080 9716 5132 9722
rect 5080 9658 5132 9664
rect 4986 9616 5042 9625
rect 4252 9580 4304 9586
rect 5814 9616 5870 9625
rect 4304 9540 4476 9568
rect 4986 9551 4988 9560
rect 4252 9522 4304 9528
rect 4160 9444 4212 9450
rect 4160 9386 4212 9392
rect 4068 9376 4120 9382
rect 4068 9318 4120 9324
rect 4055 9276 4363 9285
rect 4055 9274 4061 9276
rect 4117 9274 4141 9276
rect 4197 9274 4221 9276
rect 4277 9274 4301 9276
rect 4357 9274 4363 9276
rect 4117 9222 4119 9274
rect 4299 9222 4301 9274
rect 4055 9220 4061 9222
rect 4117 9220 4141 9222
rect 4197 9220 4221 9222
rect 4277 9220 4301 9222
rect 4357 9220 4363 9222
rect 4055 9211 4363 9220
rect 3976 9104 4028 9110
rect 3976 9046 4028 9052
rect 4160 8968 4212 8974
rect 3804 8906 3924 8922
rect 4448 8956 4476 9540
rect 5040 9551 5042 9560
rect 5172 9580 5224 9586
rect 4988 9522 5040 9528
rect 5172 9522 5224 9528
rect 5356 9580 5408 9586
rect 5356 9522 5408 9528
rect 5724 9580 5776 9586
rect 5776 9560 5814 9568
rect 5776 9551 5870 9560
rect 5776 9540 5856 9551
rect 5724 9522 5776 9528
rect 4620 9512 4672 9518
rect 4620 9454 4672 9460
rect 4896 9512 4948 9518
rect 4896 9454 4948 9460
rect 4632 9330 4660 9454
rect 4632 9302 4752 9330
rect 4724 9178 4752 9302
rect 4908 9178 4936 9454
rect 4712 9172 4764 9178
rect 4712 9114 4764 9120
rect 4896 9172 4948 9178
rect 4896 9114 4948 9120
rect 5000 9110 5028 9522
rect 5080 9376 5132 9382
rect 5080 9318 5132 9324
rect 4988 9104 5040 9110
rect 4988 9046 5040 9052
rect 4212 8928 4660 8956
rect 4160 8910 4212 8916
rect 3700 8900 3752 8906
rect 3804 8900 3936 8906
rect 3804 8894 3884 8900
rect 3700 8842 3752 8848
rect 3884 8842 3936 8848
rect 3712 8634 3740 8842
rect 3700 8628 3752 8634
rect 3700 8570 3752 8576
rect 3896 8566 3924 8842
rect 3884 8560 3936 8566
rect 3884 8502 3936 8508
rect 4436 8492 4488 8498
rect 4436 8434 4488 8440
rect 3516 8424 3568 8430
rect 3516 8366 3568 8372
rect 3240 8288 3292 8294
rect 3240 8230 3292 8236
rect 3252 7342 3280 8230
rect 3528 7410 3556 8366
rect 4055 8188 4363 8197
rect 4055 8186 4061 8188
rect 4117 8186 4141 8188
rect 4197 8186 4221 8188
rect 4277 8186 4301 8188
rect 4357 8186 4363 8188
rect 4117 8134 4119 8186
rect 4299 8134 4301 8186
rect 4055 8132 4061 8134
rect 4117 8132 4141 8134
rect 4197 8132 4221 8134
rect 4277 8132 4301 8134
rect 4357 8132 4363 8134
rect 4055 8123 4363 8132
rect 4448 7954 4476 8434
rect 4528 8356 4580 8362
rect 4528 8298 4580 8304
rect 4436 7948 4488 7954
rect 4436 7890 4488 7896
rect 3516 7404 3568 7410
rect 3516 7346 3568 7352
rect 3240 7336 3292 7342
rect 3240 7278 3292 7284
rect 3240 6384 3292 6390
rect 3240 6326 3292 6332
rect 3148 5704 3200 5710
rect 3148 5646 3200 5652
rect 2976 5358 3096 5386
rect 2872 5228 2924 5234
rect 2872 5170 2924 5176
rect 2884 4826 2912 5170
rect 2872 4820 2924 4826
rect 2872 4762 2924 4768
rect 2976 4758 3004 5358
rect 3056 5024 3108 5030
rect 3056 4966 3108 4972
rect 2964 4752 3016 4758
rect 2964 4694 3016 4700
rect 2596 4684 2648 4690
rect 2516 4644 2596 4672
rect 2596 4626 2648 4632
rect 3068 4622 3096 4966
rect 3056 4616 3108 4622
rect 3056 4558 3108 4564
rect 2645 4380 2953 4389
rect 2645 4378 2651 4380
rect 2707 4378 2731 4380
rect 2787 4378 2811 4380
rect 2867 4378 2891 4380
rect 2947 4378 2953 4380
rect 2707 4326 2709 4378
rect 2889 4326 2891 4378
rect 2645 4324 2651 4326
rect 2707 4324 2731 4326
rect 2787 4324 2811 4326
rect 2867 4324 2891 4326
rect 2947 4324 2953 4326
rect 2645 4315 2953 4324
rect 2412 3596 2464 3602
rect 2412 3538 2464 3544
rect 3252 3534 3280 6326
rect 3424 6112 3476 6118
rect 3424 6054 3476 6060
rect 3436 5914 3464 6054
rect 3424 5908 3476 5914
rect 3424 5850 3476 5856
rect 3424 5092 3476 5098
rect 3424 5034 3476 5040
rect 3436 4146 3464 5034
rect 3424 4140 3476 4146
rect 3424 4082 3476 4088
rect 3424 3936 3476 3942
rect 3424 3878 3476 3884
rect 3240 3528 3292 3534
rect 3240 3470 3292 3476
rect 3148 3460 3200 3466
rect 3148 3402 3200 3408
rect 3056 3392 3108 3398
rect 3056 3334 3108 3340
rect 2645 3292 2953 3301
rect 2645 3290 2651 3292
rect 2707 3290 2731 3292
rect 2787 3290 2811 3292
rect 2867 3290 2891 3292
rect 2947 3290 2953 3292
rect 2707 3238 2709 3290
rect 2889 3238 2891 3290
rect 2645 3236 2651 3238
rect 2707 3236 2731 3238
rect 2787 3236 2811 3238
rect 2867 3236 2891 3238
rect 2947 3236 2953 3238
rect 2645 3227 2953 3236
rect 3068 3126 3096 3334
rect 3160 3194 3188 3402
rect 3148 3188 3200 3194
rect 3148 3130 3200 3136
rect 3056 3120 3108 3126
rect 3056 3062 3108 3068
rect 2320 3052 2372 3058
rect 2320 2994 2372 3000
rect 3056 2984 3108 2990
rect 3252 2938 3280 3470
rect 3332 3460 3384 3466
rect 3332 3402 3384 3408
rect 3344 3194 3372 3402
rect 3436 3194 3464 3878
rect 3332 3188 3384 3194
rect 3332 3130 3384 3136
rect 3424 3188 3476 3194
rect 3424 3130 3476 3136
rect 3108 2932 3280 2938
rect 3056 2926 3280 2932
rect 3068 2910 3280 2926
rect 2136 2848 2188 2854
rect 2136 2790 2188 2796
rect 1985 2748 2293 2757
rect 1985 2746 1991 2748
rect 2047 2746 2071 2748
rect 2127 2746 2151 2748
rect 2207 2746 2231 2748
rect 2287 2746 2293 2748
rect 2047 2694 2049 2746
rect 2229 2694 2231 2746
rect 1985 2692 1991 2694
rect 2047 2692 2071 2694
rect 2127 2692 2151 2694
rect 2207 2692 2231 2694
rect 2287 2692 2293 2694
rect 1985 2683 2293 2692
rect 3528 2650 3556 7346
rect 4055 7100 4363 7109
rect 4055 7098 4061 7100
rect 4117 7098 4141 7100
rect 4197 7098 4221 7100
rect 4277 7098 4301 7100
rect 4357 7098 4363 7100
rect 4117 7046 4119 7098
rect 4299 7046 4301 7098
rect 4055 7044 4061 7046
rect 4117 7044 4141 7046
rect 4197 7044 4221 7046
rect 4277 7044 4301 7046
rect 4357 7044 4363 7046
rect 4055 7035 4363 7044
rect 4160 6860 4212 6866
rect 4160 6802 4212 6808
rect 3884 6724 3936 6730
rect 3884 6666 3936 6672
rect 3896 5710 3924 6666
rect 3976 6656 4028 6662
rect 3976 6598 4028 6604
rect 3988 6390 4016 6598
rect 3976 6384 4028 6390
rect 3976 6326 4028 6332
rect 4172 6322 4200 6802
rect 4540 6798 4568 8298
rect 4632 6866 4660 8928
rect 4715 8732 5023 8741
rect 4715 8730 4721 8732
rect 4777 8730 4801 8732
rect 4857 8730 4881 8732
rect 4937 8730 4961 8732
rect 5017 8730 5023 8732
rect 4777 8678 4779 8730
rect 4959 8678 4961 8730
rect 4715 8676 4721 8678
rect 4777 8676 4801 8678
rect 4857 8676 4881 8678
rect 4937 8676 4961 8678
rect 5017 8676 5023 8678
rect 4715 8667 5023 8676
rect 5092 8090 5120 9318
rect 5184 8838 5212 9522
rect 5264 9512 5316 9518
rect 5264 9454 5316 9460
rect 5276 8974 5304 9454
rect 5264 8968 5316 8974
rect 5264 8910 5316 8916
rect 5172 8832 5224 8838
rect 5172 8774 5224 8780
rect 5184 8634 5212 8774
rect 5368 8634 5396 9522
rect 5816 9376 5868 9382
rect 5816 9318 5868 9324
rect 5908 9376 5960 9382
rect 5908 9318 5960 9324
rect 6000 9376 6052 9382
rect 6000 9318 6052 9324
rect 5828 9178 5856 9318
rect 5540 9172 5592 9178
rect 5540 9114 5592 9120
rect 5816 9172 5868 9178
rect 5816 9114 5868 9120
rect 5448 8968 5500 8974
rect 5448 8910 5500 8916
rect 5172 8628 5224 8634
rect 5172 8570 5224 8576
rect 5356 8628 5408 8634
rect 5356 8570 5408 8576
rect 5080 8084 5132 8090
rect 5080 8026 5132 8032
rect 5184 7886 5212 8570
rect 5264 8492 5316 8498
rect 5264 8434 5316 8440
rect 5356 8492 5408 8498
rect 5356 8434 5408 8440
rect 5276 8022 5304 8434
rect 5264 8016 5316 8022
rect 5264 7958 5316 7964
rect 5276 7886 5304 7958
rect 5172 7880 5224 7886
rect 5172 7822 5224 7828
rect 5264 7880 5316 7886
rect 5264 7822 5316 7828
rect 5184 7750 5212 7822
rect 5172 7744 5224 7750
rect 5172 7686 5224 7692
rect 4715 7644 5023 7653
rect 4715 7642 4721 7644
rect 4777 7642 4801 7644
rect 4857 7642 4881 7644
rect 4937 7642 4961 7644
rect 5017 7642 5023 7644
rect 4777 7590 4779 7642
rect 4959 7590 4961 7642
rect 4715 7588 4721 7590
rect 4777 7588 4801 7590
rect 4857 7588 4881 7590
rect 4937 7588 4961 7590
rect 5017 7588 5023 7590
rect 4715 7579 5023 7588
rect 5172 7200 5224 7206
rect 5172 7142 5224 7148
rect 4712 6996 4764 7002
rect 4712 6938 4764 6944
rect 4620 6860 4672 6866
rect 4620 6802 4672 6808
rect 4528 6792 4580 6798
rect 4528 6734 4580 6740
rect 4344 6656 4396 6662
rect 4344 6598 4396 6604
rect 4356 6458 4384 6598
rect 4344 6452 4396 6458
rect 4344 6394 4396 6400
rect 4160 6316 4212 6322
rect 4160 6258 4212 6264
rect 4356 6254 4384 6394
rect 4344 6248 4396 6254
rect 4344 6190 4396 6196
rect 4540 6118 4568 6734
rect 4724 6644 4752 6938
rect 4632 6616 4752 6644
rect 4528 6112 4580 6118
rect 4528 6054 4580 6060
rect 4055 6012 4363 6021
rect 4055 6010 4061 6012
rect 4117 6010 4141 6012
rect 4197 6010 4221 6012
rect 4277 6010 4301 6012
rect 4357 6010 4363 6012
rect 4117 5958 4119 6010
rect 4299 5958 4301 6010
rect 4055 5956 4061 5958
rect 4117 5956 4141 5958
rect 4197 5956 4221 5958
rect 4277 5956 4301 5958
rect 4357 5956 4363 5958
rect 4055 5947 4363 5956
rect 3884 5704 3936 5710
rect 3884 5646 3936 5652
rect 4068 5704 4120 5710
rect 4068 5646 4120 5652
rect 4436 5704 4488 5710
rect 4436 5646 4488 5652
rect 3896 4622 3924 5646
rect 4080 5098 4108 5646
rect 4448 5234 4476 5646
rect 4528 5568 4580 5574
rect 4528 5510 4580 5516
rect 4436 5228 4488 5234
rect 4436 5170 4488 5176
rect 4068 5092 4120 5098
rect 4068 5034 4120 5040
rect 4055 4924 4363 4933
rect 4055 4922 4061 4924
rect 4117 4922 4141 4924
rect 4197 4922 4221 4924
rect 4277 4922 4301 4924
rect 4357 4922 4363 4924
rect 4117 4870 4119 4922
rect 4299 4870 4301 4922
rect 4055 4868 4061 4870
rect 4117 4868 4141 4870
rect 4197 4868 4221 4870
rect 4277 4868 4301 4870
rect 4357 4868 4363 4870
rect 4055 4859 4363 4868
rect 3884 4616 3936 4622
rect 3884 4558 3936 4564
rect 4068 4616 4120 4622
rect 4068 4558 4120 4564
rect 3792 4480 3844 4486
rect 3792 4422 3844 4428
rect 3804 4146 3832 4422
rect 4080 4162 4108 4558
rect 3792 4140 3844 4146
rect 3792 4082 3844 4088
rect 3988 4134 4108 4162
rect 4448 4146 4476 5170
rect 4540 5166 4568 5510
rect 4528 5160 4580 5166
rect 4528 5102 4580 5108
rect 4436 4140 4488 4146
rect 3988 4078 4016 4134
rect 4436 4082 4488 4088
rect 3976 4072 4028 4078
rect 3976 4014 4028 4020
rect 3988 3738 4016 4014
rect 4055 3836 4363 3845
rect 4055 3834 4061 3836
rect 4117 3834 4141 3836
rect 4197 3834 4221 3836
rect 4277 3834 4301 3836
rect 4357 3834 4363 3836
rect 4117 3782 4119 3834
rect 4299 3782 4301 3834
rect 4055 3780 4061 3782
rect 4117 3780 4141 3782
rect 4197 3780 4221 3782
rect 4277 3780 4301 3782
rect 4357 3780 4363 3782
rect 4055 3771 4363 3780
rect 3976 3732 4028 3738
rect 3976 3674 4028 3680
rect 4344 3664 4396 3670
rect 4344 3606 4396 3612
rect 4356 3194 4384 3606
rect 4632 3534 4660 6616
rect 4715 6556 5023 6565
rect 4715 6554 4721 6556
rect 4777 6554 4801 6556
rect 4857 6554 4881 6556
rect 4937 6554 4961 6556
rect 5017 6554 5023 6556
rect 4777 6502 4779 6554
rect 4959 6502 4961 6554
rect 4715 6500 4721 6502
rect 4777 6500 4801 6502
rect 4857 6500 4881 6502
rect 4937 6500 4961 6502
rect 5017 6500 5023 6502
rect 4715 6491 5023 6500
rect 5080 6112 5132 6118
rect 5080 6054 5132 6060
rect 5092 5710 5120 6054
rect 5080 5704 5132 5710
rect 5080 5646 5132 5652
rect 4715 5468 5023 5477
rect 4715 5466 4721 5468
rect 4777 5466 4801 5468
rect 4857 5466 4881 5468
rect 4937 5466 4961 5468
rect 5017 5466 5023 5468
rect 4777 5414 4779 5466
rect 4959 5414 4961 5466
rect 4715 5412 4721 5414
rect 4777 5412 4801 5414
rect 4857 5412 4881 5414
rect 4937 5412 4961 5414
rect 5017 5412 5023 5414
rect 4715 5403 5023 5412
rect 5092 5370 5120 5646
rect 5080 5364 5132 5370
rect 5080 5306 5132 5312
rect 5184 5098 5212 7142
rect 5276 6730 5304 7822
rect 5368 7546 5396 8434
rect 5460 8090 5488 8910
rect 5448 8084 5500 8090
rect 5448 8026 5500 8032
rect 5448 7948 5500 7954
rect 5448 7890 5500 7896
rect 5460 7546 5488 7890
rect 5356 7540 5408 7546
rect 5356 7482 5408 7488
rect 5448 7540 5500 7546
rect 5448 7482 5500 7488
rect 5552 7274 5580 9114
rect 5920 8294 5948 9318
rect 6012 8838 6040 9318
rect 6125 9276 6433 9285
rect 6125 9274 6131 9276
rect 6187 9274 6211 9276
rect 6267 9274 6291 9276
rect 6347 9274 6371 9276
rect 6427 9274 6433 9276
rect 6187 9222 6189 9274
rect 6369 9222 6371 9274
rect 6125 9220 6131 9222
rect 6187 9220 6211 9222
rect 6267 9220 6291 9222
rect 6347 9220 6371 9222
rect 6427 9220 6433 9222
rect 6125 9211 6433 9220
rect 6000 8832 6052 8838
rect 6000 8774 6052 8780
rect 6000 8356 6052 8362
rect 6000 8298 6052 8304
rect 5908 8288 5960 8294
rect 5908 8230 5960 8236
rect 5920 7954 5948 8230
rect 6012 7954 6040 8298
rect 6125 8188 6433 8197
rect 6125 8186 6131 8188
rect 6187 8186 6211 8188
rect 6267 8186 6291 8188
rect 6347 8186 6371 8188
rect 6427 8186 6433 8188
rect 6187 8134 6189 8186
rect 6369 8134 6371 8186
rect 6125 8132 6131 8134
rect 6187 8132 6211 8134
rect 6267 8132 6291 8134
rect 6347 8132 6371 8134
rect 6427 8132 6433 8134
rect 6125 8123 6433 8132
rect 5908 7948 5960 7954
rect 5908 7890 5960 7896
rect 6000 7948 6052 7954
rect 6000 7890 6052 7896
rect 5908 7744 5960 7750
rect 5908 7686 5960 7692
rect 5540 7268 5592 7274
rect 5540 7210 5592 7216
rect 5264 6724 5316 6730
rect 5264 6666 5316 6672
rect 5356 5908 5408 5914
rect 5356 5850 5408 5856
rect 5368 5234 5396 5850
rect 5816 5636 5868 5642
rect 5816 5578 5868 5584
rect 5356 5228 5408 5234
rect 5356 5170 5408 5176
rect 5632 5228 5684 5234
rect 5632 5170 5684 5176
rect 5172 5092 5224 5098
rect 5172 5034 5224 5040
rect 4896 5024 4948 5030
rect 4896 4966 4948 4972
rect 4908 4826 4936 4966
rect 4896 4820 4948 4826
rect 4896 4762 4948 4768
rect 5080 4616 5132 4622
rect 5080 4558 5132 4564
rect 4715 4380 5023 4389
rect 4715 4378 4721 4380
rect 4777 4378 4801 4380
rect 4857 4378 4881 4380
rect 4937 4378 4961 4380
rect 5017 4378 5023 4380
rect 4777 4326 4779 4378
rect 4959 4326 4961 4378
rect 4715 4324 4721 4326
rect 4777 4324 4801 4326
rect 4857 4324 4881 4326
rect 4937 4324 4961 4326
rect 5017 4324 5023 4326
rect 4715 4315 5023 4324
rect 5092 3738 5120 4558
rect 5184 4486 5212 5034
rect 5368 4554 5396 5170
rect 5448 5024 5500 5030
rect 5448 4966 5500 4972
rect 5460 4826 5488 4966
rect 5448 4820 5500 4826
rect 5448 4762 5500 4768
rect 5540 4752 5592 4758
rect 5540 4694 5592 4700
rect 5356 4548 5408 4554
rect 5356 4490 5408 4496
rect 5172 4480 5224 4486
rect 5172 4422 5224 4428
rect 5552 3738 5580 4694
rect 5644 4486 5672 5170
rect 5632 4480 5684 4486
rect 5632 4422 5684 4428
rect 5724 4480 5776 4486
rect 5724 4422 5776 4428
rect 5080 3732 5132 3738
rect 5080 3674 5132 3680
rect 5540 3732 5592 3738
rect 5540 3674 5592 3680
rect 5552 3618 5580 3674
rect 5460 3590 5580 3618
rect 4436 3528 4488 3534
rect 4436 3470 4488 3476
rect 4620 3528 4672 3534
rect 4620 3470 4672 3476
rect 5356 3528 5408 3534
rect 5356 3470 5408 3476
rect 4448 3194 4476 3470
rect 4344 3188 4396 3194
rect 4344 3130 4396 3136
rect 4436 3188 4488 3194
rect 4436 3130 4488 3136
rect 4632 3058 4660 3470
rect 5080 3392 5132 3398
rect 5080 3334 5132 3340
rect 4715 3292 5023 3301
rect 4715 3290 4721 3292
rect 4777 3290 4801 3292
rect 4857 3290 4881 3292
rect 4937 3290 4961 3292
rect 5017 3290 5023 3292
rect 4777 3238 4779 3290
rect 4959 3238 4961 3290
rect 4715 3236 4721 3238
rect 4777 3236 4801 3238
rect 4857 3236 4881 3238
rect 4937 3236 4961 3238
rect 5017 3236 5023 3238
rect 4715 3227 5023 3236
rect 5092 3058 5120 3334
rect 4620 3052 4672 3058
rect 4620 2994 4672 3000
rect 5080 3052 5132 3058
rect 5080 2994 5132 3000
rect 4436 2984 4488 2990
rect 4436 2926 4488 2932
rect 4055 2748 4363 2757
rect 4055 2746 4061 2748
rect 4117 2746 4141 2748
rect 4197 2746 4221 2748
rect 4277 2746 4301 2748
rect 4357 2746 4363 2748
rect 4117 2694 4119 2746
rect 4299 2694 4301 2746
rect 4055 2692 4061 2694
rect 4117 2692 4141 2694
rect 4197 2692 4221 2694
rect 4277 2692 4301 2694
rect 4357 2692 4363 2694
rect 4055 2683 4363 2692
rect 4448 2650 4476 2926
rect 5368 2922 5396 3470
rect 5460 3058 5488 3590
rect 5540 3528 5592 3534
rect 5540 3470 5592 3476
rect 5552 3194 5580 3470
rect 5540 3188 5592 3194
rect 5540 3130 5592 3136
rect 5448 3052 5500 3058
rect 5632 3052 5684 3058
rect 5500 3012 5580 3040
rect 5448 2994 5500 3000
rect 5356 2916 5408 2922
rect 5356 2858 5408 2864
rect 5368 2774 5396 2858
rect 5368 2746 5488 2774
rect 3516 2644 3568 2650
rect 3516 2586 3568 2592
rect 4436 2644 4488 2650
rect 4436 2586 4488 2592
rect 1308 2508 1360 2514
rect 1308 2450 1360 2456
rect 1216 2440 1268 2446
rect 1216 2382 1268 2388
rect 20 2372 72 2378
rect 20 2314 72 2320
rect 32 800 60 2314
rect 1228 1465 1256 2382
rect 1214 1456 1270 1465
rect 1214 1391 1270 1400
rect 1320 800 1348 2450
rect 5460 2446 5488 2746
rect 5552 2446 5580 3012
rect 5632 2994 5684 3000
rect 5644 2650 5672 2994
rect 5736 2854 5764 4422
rect 5724 2848 5776 2854
rect 5724 2790 5776 2796
rect 5632 2644 5684 2650
rect 5632 2586 5684 2592
rect 5828 2446 5856 5578
rect 5920 2774 5948 7686
rect 6012 7546 6040 7890
rect 6368 7880 6420 7886
rect 6368 7822 6420 7828
rect 6092 7812 6144 7818
rect 6092 7754 6144 7760
rect 6000 7540 6052 7546
rect 6000 7482 6052 7488
rect 6104 7188 6132 7754
rect 6380 7342 6408 7822
rect 6368 7336 6420 7342
rect 6368 7278 6420 7284
rect 6012 7160 6132 7188
rect 6012 7002 6040 7160
rect 6125 7100 6433 7109
rect 6125 7098 6131 7100
rect 6187 7098 6211 7100
rect 6267 7098 6291 7100
rect 6347 7098 6371 7100
rect 6427 7098 6433 7100
rect 6187 7046 6189 7098
rect 6369 7046 6371 7098
rect 6125 7044 6131 7046
rect 6187 7044 6211 7046
rect 6267 7044 6291 7046
rect 6347 7044 6371 7046
rect 6427 7044 6433 7046
rect 6125 7035 6433 7044
rect 6000 6996 6052 7002
rect 6000 6938 6052 6944
rect 6012 6458 6040 6938
rect 6656 6798 6684 9862
rect 6785 9820 7093 9829
rect 6785 9818 6791 9820
rect 6847 9818 6871 9820
rect 6927 9818 6951 9820
rect 7007 9818 7031 9820
rect 7087 9818 7093 9820
rect 6847 9766 6849 9818
rect 7029 9766 7031 9818
rect 6785 9764 6791 9766
rect 6847 9764 6871 9766
rect 6927 9764 6951 9766
rect 7007 9764 7031 9766
rect 7087 9764 7093 9766
rect 6785 9755 7093 9764
rect 6920 9580 6972 9586
rect 6920 9522 6972 9528
rect 6932 9110 6960 9522
rect 6920 9104 6972 9110
rect 6920 9046 6972 9052
rect 6932 8974 6960 9046
rect 6920 8968 6972 8974
rect 6920 8910 6972 8916
rect 6785 8732 7093 8741
rect 6785 8730 6791 8732
rect 6847 8730 6871 8732
rect 6927 8730 6951 8732
rect 7007 8730 7031 8732
rect 7087 8730 7093 8732
rect 6847 8678 6849 8730
rect 7029 8678 7031 8730
rect 6785 8676 6791 8678
rect 6847 8676 6871 8678
rect 6927 8676 6951 8678
rect 7007 8676 7031 8678
rect 7087 8676 7093 8678
rect 6785 8667 7093 8676
rect 6920 8628 6972 8634
rect 6920 8570 6972 8576
rect 6932 8090 6960 8570
rect 7012 8492 7064 8498
rect 7012 8434 7064 8440
rect 7196 8492 7248 8498
rect 7196 8434 7248 8440
rect 6920 8084 6972 8090
rect 6920 8026 6972 8032
rect 7024 7750 7052 8434
rect 7208 8090 7236 8434
rect 7196 8084 7248 8090
rect 7196 8026 7248 8032
rect 7196 7880 7248 7886
rect 7196 7822 7248 7828
rect 7012 7744 7064 7750
rect 7012 7686 7064 7692
rect 6785 7644 7093 7653
rect 6785 7642 6791 7644
rect 6847 7642 6871 7644
rect 6927 7642 6951 7644
rect 7007 7642 7031 7644
rect 7087 7642 7093 7644
rect 6847 7590 6849 7642
rect 7029 7590 7031 7642
rect 6785 7588 6791 7590
rect 6847 7588 6871 7590
rect 6927 7588 6951 7590
rect 7007 7588 7031 7590
rect 7087 7588 7093 7590
rect 6785 7579 7093 7588
rect 7208 7342 7236 7822
rect 7196 7336 7248 7342
rect 7196 7278 7248 7284
rect 6644 6792 6696 6798
rect 6644 6734 6696 6740
rect 7196 6792 7248 6798
rect 7196 6734 7248 6740
rect 6000 6452 6052 6458
rect 6000 6394 6052 6400
rect 6656 6390 6684 6734
rect 6785 6556 7093 6565
rect 6785 6554 6791 6556
rect 6847 6554 6871 6556
rect 6927 6554 6951 6556
rect 7007 6554 7031 6556
rect 7087 6554 7093 6556
rect 6847 6502 6849 6554
rect 7029 6502 7031 6554
rect 6785 6500 6791 6502
rect 6847 6500 6871 6502
rect 6927 6500 6951 6502
rect 7007 6500 7031 6502
rect 7087 6500 7093 6502
rect 6785 6491 7093 6500
rect 6644 6384 6696 6390
rect 6644 6326 6696 6332
rect 6125 6012 6433 6021
rect 6125 6010 6131 6012
rect 6187 6010 6211 6012
rect 6267 6010 6291 6012
rect 6347 6010 6371 6012
rect 6427 6010 6433 6012
rect 6187 5958 6189 6010
rect 6369 5958 6371 6010
rect 6125 5956 6131 5958
rect 6187 5956 6211 5958
rect 6267 5956 6291 5958
rect 6347 5956 6371 5958
rect 6427 5956 6433 5958
rect 6125 5947 6433 5956
rect 6656 5914 6684 6326
rect 6828 6112 6880 6118
rect 6828 6054 6880 6060
rect 6644 5908 6696 5914
rect 6644 5850 6696 5856
rect 6840 5556 6868 6054
rect 7208 5914 7236 6734
rect 7196 5908 7248 5914
rect 7196 5850 7248 5856
rect 6472 5528 6868 5556
rect 6125 4924 6433 4933
rect 6125 4922 6131 4924
rect 6187 4922 6211 4924
rect 6267 4922 6291 4924
rect 6347 4922 6371 4924
rect 6427 4922 6433 4924
rect 6187 4870 6189 4922
rect 6369 4870 6371 4922
rect 6125 4868 6131 4870
rect 6187 4868 6211 4870
rect 6267 4868 6291 4870
rect 6347 4868 6371 4870
rect 6427 4868 6433 4870
rect 6125 4859 6433 4868
rect 6125 3836 6433 3845
rect 6125 3834 6131 3836
rect 6187 3834 6211 3836
rect 6267 3834 6291 3836
rect 6347 3834 6371 3836
rect 6427 3834 6433 3836
rect 6187 3782 6189 3834
rect 6369 3782 6371 3834
rect 6125 3780 6131 3782
rect 6187 3780 6211 3782
rect 6267 3780 6291 3782
rect 6347 3780 6371 3782
rect 6427 3780 6433 3782
rect 6125 3771 6433 3780
rect 6472 3058 6500 5528
rect 6785 5468 7093 5477
rect 6785 5466 6791 5468
rect 6847 5466 6871 5468
rect 6927 5466 6951 5468
rect 7007 5466 7031 5468
rect 7087 5466 7093 5468
rect 6847 5414 6849 5466
rect 7029 5414 7031 5466
rect 6785 5412 6791 5414
rect 6847 5412 6871 5414
rect 6927 5412 6951 5414
rect 7007 5412 7031 5414
rect 7087 5412 7093 5414
rect 6785 5403 7093 5412
rect 7300 5114 7328 9930
rect 7932 9920 7984 9926
rect 7932 9862 7984 9868
rect 8392 9920 8444 9926
rect 8392 9862 8444 9868
rect 7378 9616 7434 9625
rect 7434 9560 7512 9568
rect 7378 9551 7380 9560
rect 7432 9540 7512 9560
rect 7380 9522 7432 9528
rect 7380 8084 7432 8090
rect 7380 8026 7432 8032
rect 7392 7886 7420 8026
rect 7380 7880 7432 7886
rect 7380 7822 7432 7828
rect 7380 6928 7432 6934
rect 7380 6870 7432 6876
rect 7116 5086 7328 5114
rect 6552 5024 6604 5030
rect 6552 4966 6604 4972
rect 6564 4146 6592 4966
rect 7116 4826 7144 5086
rect 7196 5024 7248 5030
rect 7196 4966 7248 4972
rect 7208 4826 7236 4966
rect 7104 4820 7156 4826
rect 7104 4762 7156 4768
rect 7196 4820 7248 4826
rect 7196 4762 7248 4768
rect 7288 4684 7340 4690
rect 7288 4626 7340 4632
rect 6644 4616 6696 4622
rect 6644 4558 6696 4564
rect 6552 4140 6604 4146
rect 6552 4082 6604 4088
rect 6460 3052 6512 3058
rect 6460 2994 6512 3000
rect 5920 2746 6040 2774
rect 6012 2650 6040 2746
rect 6125 2748 6433 2757
rect 6125 2746 6131 2748
rect 6187 2746 6211 2748
rect 6267 2746 6291 2748
rect 6347 2746 6371 2748
rect 6427 2746 6433 2748
rect 6187 2694 6189 2746
rect 6369 2694 6371 2746
rect 6125 2692 6131 2694
rect 6187 2692 6211 2694
rect 6267 2692 6291 2694
rect 6347 2692 6371 2694
rect 6427 2692 6433 2694
rect 6125 2683 6433 2692
rect 6656 2650 6684 4558
rect 7196 4480 7248 4486
rect 7196 4422 7248 4428
rect 6785 4380 7093 4389
rect 6785 4378 6791 4380
rect 6847 4378 6871 4380
rect 6927 4378 6951 4380
rect 7007 4378 7031 4380
rect 7087 4378 7093 4380
rect 6847 4326 6849 4378
rect 7029 4326 7031 4378
rect 6785 4324 6791 4326
rect 6847 4324 6871 4326
rect 6927 4324 6951 4326
rect 7007 4324 7031 4326
rect 7087 4324 7093 4326
rect 6785 4315 7093 4324
rect 7208 4162 7236 4422
rect 7300 4282 7328 4626
rect 7288 4276 7340 4282
rect 7288 4218 7340 4224
rect 7208 4134 7328 4162
rect 7300 4078 7328 4134
rect 7288 4072 7340 4078
rect 7288 4014 7340 4020
rect 7196 3528 7248 3534
rect 7196 3470 7248 3476
rect 6785 3292 7093 3301
rect 6785 3290 6791 3292
rect 6847 3290 6871 3292
rect 6927 3290 6951 3292
rect 7007 3290 7031 3292
rect 7087 3290 7093 3292
rect 6847 3238 6849 3290
rect 7029 3238 7031 3290
rect 6785 3236 6791 3238
rect 6847 3236 6871 3238
rect 6927 3236 6951 3238
rect 7007 3236 7031 3238
rect 7087 3236 7093 3238
rect 6785 3227 7093 3236
rect 7208 3058 7236 3470
rect 7300 3194 7328 4014
rect 7392 3942 7420 6870
rect 7484 6118 7512 9540
rect 7944 9518 7972 9862
rect 8404 9722 8432 9862
rect 8392 9716 8444 9722
rect 8392 9658 8444 9664
rect 7932 9512 7984 9518
rect 7932 9454 7984 9460
rect 8116 9512 8168 9518
rect 8116 9454 8168 9460
rect 7748 9376 7800 9382
rect 7748 9318 7800 9324
rect 7760 9042 7788 9318
rect 7840 9104 7892 9110
rect 7840 9046 7892 9052
rect 7748 9036 7800 9042
rect 7748 8978 7800 8984
rect 7564 8628 7616 8634
rect 7616 8588 7696 8616
rect 7564 8570 7616 8576
rect 7564 8288 7616 8294
rect 7564 8230 7616 8236
rect 7576 8090 7604 8230
rect 7668 8090 7696 8588
rect 7564 8084 7616 8090
rect 7564 8026 7616 8032
rect 7656 8084 7708 8090
rect 7656 8026 7708 8032
rect 7760 6934 7788 8978
rect 7748 6928 7800 6934
rect 7748 6870 7800 6876
rect 7656 6792 7708 6798
rect 7656 6734 7708 6740
rect 7668 6458 7696 6734
rect 7852 6662 7880 9046
rect 8024 9036 8076 9042
rect 8024 8978 8076 8984
rect 7932 8968 7984 8974
rect 7932 8910 7984 8916
rect 7944 8634 7972 8910
rect 7932 8628 7984 8634
rect 7932 8570 7984 8576
rect 8036 8430 8064 8978
rect 8024 8424 8076 8430
rect 8024 8366 8076 8372
rect 8036 8090 8064 8366
rect 8024 8084 8076 8090
rect 8024 8026 8076 8032
rect 8128 7818 8156 9454
rect 8195 9276 8503 9285
rect 8195 9274 8201 9276
rect 8257 9274 8281 9276
rect 8337 9274 8361 9276
rect 8417 9274 8441 9276
rect 8497 9274 8503 9276
rect 8257 9222 8259 9274
rect 8439 9222 8441 9274
rect 8195 9220 8201 9222
rect 8257 9220 8281 9222
rect 8337 9220 8361 9222
rect 8417 9220 8441 9222
rect 8497 9220 8503 9222
rect 8195 9211 8503 9220
rect 8588 9178 8616 10016
rect 8668 9998 8720 10004
rect 8680 9518 8708 9998
rect 8760 9920 8812 9926
rect 8760 9862 8812 9868
rect 8772 9654 8800 9862
rect 8855 9820 9163 9829
rect 8855 9818 8861 9820
rect 8917 9818 8941 9820
rect 8997 9818 9021 9820
rect 9077 9818 9101 9820
rect 9157 9818 9163 9820
rect 8917 9766 8919 9818
rect 9099 9766 9101 9818
rect 8855 9764 8861 9766
rect 8917 9764 8941 9766
rect 8997 9764 9021 9766
rect 9077 9764 9101 9766
rect 9157 9764 9163 9766
rect 8855 9755 9163 9764
rect 8760 9648 8812 9654
rect 8760 9590 8812 9596
rect 8668 9512 8720 9518
rect 8668 9454 8720 9460
rect 8576 9172 8628 9178
rect 8576 9114 8628 9120
rect 9324 8974 9352 11591
rect 9402 10296 9458 10305
rect 9402 10231 9458 10240
rect 9416 9722 9444 10231
rect 9692 10062 9720 11911
rect 9680 10056 9732 10062
rect 9680 9998 9732 10004
rect 9404 9716 9456 9722
rect 9404 9658 9456 9664
rect 9312 8968 9364 8974
rect 9312 8910 9364 8916
rect 8855 8732 9163 8741
rect 8855 8730 8861 8732
rect 8917 8730 8941 8732
rect 8997 8730 9021 8732
rect 9077 8730 9101 8732
rect 9157 8730 9163 8732
rect 8917 8678 8919 8730
rect 9099 8678 9101 8730
rect 8855 8676 8861 8678
rect 8917 8676 8941 8678
rect 8997 8676 9021 8678
rect 9077 8676 9101 8678
rect 9157 8676 9163 8678
rect 8855 8667 9163 8676
rect 8668 8492 8720 8498
rect 8668 8434 8720 8440
rect 8195 8188 8503 8197
rect 8195 8186 8201 8188
rect 8257 8186 8281 8188
rect 8337 8186 8361 8188
rect 8417 8186 8441 8188
rect 8497 8186 8503 8188
rect 8257 8134 8259 8186
rect 8439 8134 8441 8186
rect 8195 8132 8201 8134
rect 8257 8132 8281 8134
rect 8337 8132 8361 8134
rect 8417 8132 8441 8134
rect 8497 8132 8503 8134
rect 8195 8123 8503 8132
rect 8576 8084 8628 8090
rect 8576 8026 8628 8032
rect 8116 7812 8168 7818
rect 8116 7754 8168 7760
rect 8024 7268 8076 7274
rect 8024 7210 8076 7216
rect 8036 6934 8064 7210
rect 8024 6928 8076 6934
rect 8024 6870 8076 6876
rect 7932 6792 7984 6798
rect 7932 6734 7984 6740
rect 7840 6656 7892 6662
rect 7840 6598 7892 6604
rect 7656 6452 7708 6458
rect 7656 6394 7708 6400
rect 7668 6322 7696 6394
rect 7564 6316 7616 6322
rect 7564 6258 7616 6264
rect 7656 6316 7708 6322
rect 7656 6258 7708 6264
rect 7576 6118 7604 6258
rect 7472 6112 7524 6118
rect 7472 6054 7524 6060
rect 7564 6112 7616 6118
rect 7564 6054 7616 6060
rect 7656 6112 7708 6118
rect 7656 6054 7708 6060
rect 7576 5642 7604 6054
rect 7668 5710 7696 6054
rect 7852 5794 7880 6598
rect 7944 6186 7972 6734
rect 7932 6180 7984 6186
rect 7932 6122 7984 6128
rect 7944 5914 7972 6122
rect 7932 5908 7984 5914
rect 7932 5850 7984 5856
rect 8128 5794 8156 7754
rect 8484 7744 8536 7750
rect 8484 7686 8536 7692
rect 8496 7274 8524 7686
rect 8588 7342 8616 8026
rect 8680 7546 8708 8434
rect 9036 8356 9088 8362
rect 9036 8298 9088 8304
rect 9048 8265 9076 8298
rect 9034 8256 9090 8265
rect 9034 8191 9090 8200
rect 8855 7644 9163 7653
rect 8855 7642 8861 7644
rect 8917 7642 8941 7644
rect 8997 7642 9021 7644
rect 9077 7642 9101 7644
rect 9157 7642 9163 7644
rect 8917 7590 8919 7642
rect 9099 7590 9101 7642
rect 8855 7588 8861 7590
rect 8917 7588 8941 7590
rect 8997 7588 9021 7590
rect 9077 7588 9101 7590
rect 9157 7588 9163 7590
rect 8855 7579 9163 7588
rect 8668 7540 8720 7546
rect 8668 7482 8720 7488
rect 8668 7404 8720 7410
rect 8668 7346 8720 7352
rect 8576 7336 8628 7342
rect 8576 7278 8628 7284
rect 8484 7268 8536 7274
rect 8484 7210 8536 7216
rect 8195 7100 8503 7109
rect 8195 7098 8201 7100
rect 8257 7098 8281 7100
rect 8337 7098 8361 7100
rect 8417 7098 8441 7100
rect 8497 7098 8503 7100
rect 8257 7046 8259 7098
rect 8439 7046 8441 7098
rect 8195 7044 8201 7046
rect 8257 7044 8281 7046
rect 8337 7044 8361 7046
rect 8417 7044 8441 7046
rect 8497 7044 8503 7046
rect 8195 7035 8503 7044
rect 8588 6984 8616 7278
rect 8496 6956 8616 6984
rect 8392 6792 8444 6798
rect 8392 6734 8444 6740
rect 8208 6656 8260 6662
rect 8208 6598 8260 6604
rect 8220 6458 8248 6598
rect 8208 6452 8260 6458
rect 8208 6394 8260 6400
rect 8404 6322 8432 6734
rect 8496 6662 8524 6956
rect 8484 6656 8536 6662
rect 8484 6598 8536 6604
rect 8392 6316 8444 6322
rect 8392 6258 8444 6264
rect 8496 6202 8524 6598
rect 8680 6458 8708 7346
rect 8855 6556 9163 6565
rect 8855 6554 8861 6556
rect 8917 6554 8941 6556
rect 8997 6554 9021 6556
rect 9077 6554 9101 6556
rect 9157 6554 9163 6556
rect 8917 6502 8919 6554
rect 9099 6502 9101 6554
rect 8855 6500 8861 6502
rect 8917 6500 8941 6502
rect 8997 6500 9021 6502
rect 9077 6500 9101 6502
rect 9157 6500 9163 6502
rect 8855 6491 9163 6500
rect 8668 6452 8720 6458
rect 8668 6394 8720 6400
rect 8666 6216 8722 6225
rect 8496 6186 8616 6202
rect 8484 6180 8616 6186
rect 8536 6174 8616 6180
rect 8484 6122 8536 6128
rect 8195 6012 8503 6021
rect 8195 6010 8201 6012
rect 8257 6010 8281 6012
rect 8337 6010 8361 6012
rect 8417 6010 8441 6012
rect 8497 6010 8503 6012
rect 8257 5958 8259 6010
rect 8439 5958 8441 6010
rect 8195 5956 8201 5958
rect 8257 5956 8281 5958
rect 8337 5956 8361 5958
rect 8417 5956 8441 5958
rect 8497 5956 8503 5958
rect 8195 5947 8503 5956
rect 7852 5766 7972 5794
rect 8128 5766 8248 5794
rect 7656 5704 7708 5710
rect 7656 5646 7708 5652
rect 7564 5636 7616 5642
rect 7564 5578 7616 5584
rect 7564 5160 7616 5166
rect 7564 5102 7616 5108
rect 7380 3936 7432 3942
rect 7380 3878 7432 3884
rect 7380 3596 7432 3602
rect 7380 3538 7432 3544
rect 7472 3596 7524 3602
rect 7472 3538 7524 3544
rect 7392 3194 7420 3538
rect 7288 3188 7340 3194
rect 7288 3130 7340 3136
rect 7380 3188 7432 3194
rect 7380 3130 7432 3136
rect 7196 3052 7248 3058
rect 7196 2994 7248 3000
rect 6736 2848 6788 2854
rect 6736 2790 6788 2796
rect 6000 2644 6052 2650
rect 6000 2586 6052 2592
rect 6644 2644 6696 2650
rect 6644 2586 6696 2592
rect 6748 2582 6776 2790
rect 6736 2576 6788 2582
rect 6736 2518 6788 2524
rect 7208 2514 7236 2994
rect 7380 2848 7432 2854
rect 7484 2802 7512 3538
rect 7576 3194 7604 5102
rect 7668 4758 7696 5646
rect 7748 5160 7800 5166
rect 7748 5102 7800 5108
rect 7840 5160 7892 5166
rect 7840 5102 7892 5108
rect 7656 4752 7708 4758
rect 7656 4694 7708 4700
rect 7760 4078 7788 5102
rect 7852 4826 7880 5102
rect 7840 4820 7892 4826
rect 7840 4762 7892 4768
rect 7944 4706 7972 5766
rect 8024 5704 8076 5710
rect 8024 5646 8076 5652
rect 8036 5370 8064 5646
rect 8116 5568 8168 5574
rect 8116 5510 8168 5516
rect 8024 5364 8076 5370
rect 8024 5306 8076 5312
rect 8024 5160 8076 5166
rect 8024 5102 8076 5108
rect 8036 4758 8064 5102
rect 7852 4678 7972 4706
rect 8024 4752 8076 4758
rect 8024 4694 8076 4700
rect 7748 4072 7800 4078
rect 7748 4014 7800 4020
rect 7748 3936 7800 3942
rect 7748 3878 7800 3884
rect 7760 3398 7788 3878
rect 7748 3392 7800 3398
rect 7748 3334 7800 3340
rect 7564 3188 7616 3194
rect 7564 3130 7616 3136
rect 7564 3052 7616 3058
rect 7564 2994 7616 3000
rect 7432 2796 7512 2802
rect 7380 2790 7512 2796
rect 7392 2774 7512 2790
rect 7196 2508 7248 2514
rect 7196 2450 7248 2456
rect 5448 2440 5500 2446
rect 5448 2382 5500 2388
rect 5540 2440 5592 2446
rect 5540 2382 5592 2388
rect 5816 2440 5868 2446
rect 5816 2382 5868 2388
rect 7392 2378 7420 2774
rect 7576 2650 7604 2994
rect 7760 2938 7788 3334
rect 7668 2910 7788 2938
rect 7564 2644 7616 2650
rect 7564 2586 7616 2592
rect 7564 2440 7616 2446
rect 7668 2428 7696 2910
rect 7852 2774 7880 4678
rect 8128 4622 8156 5510
rect 8220 5234 8248 5766
rect 8208 5228 8260 5234
rect 8208 5170 8260 5176
rect 8195 4924 8503 4933
rect 8195 4922 8201 4924
rect 8257 4922 8281 4924
rect 8337 4922 8361 4924
rect 8417 4922 8441 4924
rect 8497 4922 8503 4924
rect 8257 4870 8259 4922
rect 8439 4870 8441 4922
rect 8195 4868 8201 4870
rect 8257 4868 8281 4870
rect 8337 4868 8361 4870
rect 8417 4868 8441 4870
rect 8497 4868 8503 4870
rect 8195 4859 8503 4868
rect 8116 4616 8168 4622
rect 8116 4558 8168 4564
rect 8128 3058 8156 4558
rect 8195 3836 8503 3845
rect 8195 3834 8201 3836
rect 8257 3834 8281 3836
rect 8337 3834 8361 3836
rect 8417 3834 8441 3836
rect 8497 3834 8503 3836
rect 8257 3782 8259 3834
rect 8439 3782 8441 3834
rect 8195 3780 8201 3782
rect 8257 3780 8281 3782
rect 8337 3780 8361 3782
rect 8417 3780 8441 3782
rect 8497 3780 8503 3782
rect 8195 3771 8503 3780
rect 8588 3194 8616 6174
rect 8666 6151 8722 6160
rect 8680 5914 8708 6151
rect 8668 5908 8720 5914
rect 8668 5850 8720 5856
rect 8855 5468 9163 5477
rect 8855 5466 8861 5468
rect 8917 5466 8941 5468
rect 8997 5466 9021 5468
rect 9077 5466 9101 5468
rect 9157 5466 9163 5468
rect 8917 5414 8919 5466
rect 9099 5414 9101 5466
rect 8855 5412 8861 5414
rect 8917 5412 8941 5414
rect 8997 5412 9021 5414
rect 9077 5412 9101 5414
rect 9157 5412 9163 5414
rect 8855 5403 9163 5412
rect 9036 5160 9088 5166
rect 9036 5102 9088 5108
rect 9048 4865 9076 5102
rect 9034 4856 9090 4865
rect 9034 4791 9090 4800
rect 8855 4380 9163 4389
rect 8855 4378 8861 4380
rect 8917 4378 8941 4380
rect 8997 4378 9021 4380
rect 9077 4378 9101 4380
rect 9157 4378 9163 4380
rect 8917 4326 8919 4378
rect 9099 4326 9101 4378
rect 8855 4324 8861 4326
rect 8917 4324 8941 4326
rect 8997 4324 9021 4326
rect 9077 4324 9101 4326
rect 9157 4324 9163 4326
rect 8855 4315 9163 4324
rect 8668 3528 8720 3534
rect 8668 3470 8720 3476
rect 8576 3188 8628 3194
rect 8576 3130 8628 3136
rect 7932 3052 7984 3058
rect 7932 2994 7984 3000
rect 8116 3052 8168 3058
rect 8116 2994 8168 3000
rect 7944 2938 7972 2994
rect 7944 2910 8064 2938
rect 7852 2746 7972 2774
rect 7616 2400 7696 2428
rect 7564 2382 7616 2388
rect 7944 2378 7972 2746
rect 3240 2372 3292 2378
rect 3240 2314 3292 2320
rect 5724 2372 5776 2378
rect 5724 2314 5776 2320
rect 7380 2372 7432 2378
rect 7380 2314 7432 2320
rect 7748 2372 7800 2378
rect 7748 2314 7800 2320
rect 7932 2372 7984 2378
rect 7932 2314 7984 2320
rect 2645 2204 2953 2213
rect 2645 2202 2651 2204
rect 2707 2202 2731 2204
rect 2787 2202 2811 2204
rect 2867 2202 2891 2204
rect 2947 2202 2953 2204
rect 2707 2150 2709 2202
rect 2889 2150 2891 2202
rect 2645 2148 2651 2150
rect 2707 2148 2731 2150
rect 2787 2148 2811 2150
rect 2867 2148 2891 2150
rect 2947 2148 2953 2150
rect 2645 2139 2953 2148
rect 3252 800 3280 2314
rect 5632 2304 5684 2310
rect 5632 2246 5684 2252
rect 4715 2204 5023 2213
rect 4715 2202 4721 2204
rect 4777 2202 4801 2204
rect 4857 2202 4881 2204
rect 4937 2202 4961 2204
rect 5017 2202 5023 2204
rect 4777 2150 4779 2202
rect 4959 2150 4961 2202
rect 4715 2148 4721 2150
rect 4777 2148 4801 2150
rect 4857 2148 4881 2150
rect 4937 2148 4961 2150
rect 5017 2148 5023 2150
rect 4715 2139 5023 2148
rect 5644 1442 5672 2246
rect 5736 2106 5764 2314
rect 6552 2304 6604 2310
rect 6552 2246 6604 2252
rect 5724 2100 5776 2106
rect 5724 2042 5776 2048
rect 5460 1414 5672 1442
rect 5184 870 5304 898
rect 5184 800 5212 870
rect 18 0 74 800
rect 1306 0 1362 800
rect 3238 0 3294 800
rect 5170 0 5226 800
rect 5276 762 5304 870
rect 5460 762 5488 1414
rect 6564 1170 6592 2246
rect 6785 2204 7093 2213
rect 6785 2202 6791 2204
rect 6847 2202 6871 2204
rect 6927 2202 6951 2204
rect 7007 2202 7031 2204
rect 7087 2202 7093 2204
rect 6847 2150 6849 2202
rect 7029 2150 7031 2202
rect 6785 2148 6791 2150
rect 6847 2148 6871 2150
rect 6927 2148 6951 2150
rect 7007 2148 7031 2150
rect 7087 2148 7093 2150
rect 6785 2139 7093 2148
rect 7760 2106 7788 2314
rect 7748 2100 7800 2106
rect 7748 2042 7800 2048
rect 6472 1142 6592 1170
rect 6472 800 6500 1142
rect 5276 734 5488 762
rect 6458 0 6514 800
rect 8036 785 8064 2910
rect 8195 2748 8503 2757
rect 8195 2746 8201 2748
rect 8257 2746 8281 2748
rect 8337 2746 8361 2748
rect 8417 2746 8441 2748
rect 8497 2746 8503 2748
rect 8257 2694 8259 2746
rect 8439 2694 8441 2746
rect 8195 2692 8201 2694
rect 8257 2692 8281 2694
rect 8337 2692 8361 2694
rect 8417 2692 8441 2694
rect 8497 2692 8503 2694
rect 8195 2683 8503 2692
rect 8404 870 8524 898
rect 8404 800 8432 870
rect 8022 776 8078 785
rect 8022 711 8078 720
rect 8390 0 8446 800
rect 8496 762 8524 870
rect 8680 762 8708 3470
rect 8855 3292 9163 3301
rect 8855 3290 8861 3292
rect 8917 3290 8941 3292
rect 8997 3290 9021 3292
rect 9077 3290 9101 3292
rect 9157 3290 9163 3292
rect 8917 3238 8919 3290
rect 9099 3238 9101 3290
rect 8855 3236 8861 3238
rect 8917 3236 8941 3238
rect 8997 3236 9021 3238
rect 9077 3236 9101 3238
rect 9157 3236 9163 3238
rect 8855 3227 9163 3236
rect 9404 3052 9456 3058
rect 9404 2994 9456 3000
rect 9416 2825 9444 2994
rect 9402 2816 9458 2825
rect 9402 2751 9458 2760
rect 10324 2372 10376 2378
rect 10324 2314 10376 2320
rect 8855 2204 9163 2213
rect 8855 2202 8861 2204
rect 8917 2202 8941 2204
rect 8997 2202 9021 2204
rect 9077 2202 9101 2204
rect 9157 2202 9163 2204
rect 8917 2150 8919 2202
rect 9099 2150 9101 2202
rect 8855 2148 8861 2150
rect 8917 2148 8941 2150
rect 8997 2148 9021 2150
rect 9077 2148 9101 2150
rect 9157 2148 9163 2150
rect 8855 2139 9163 2148
rect 10336 800 10364 2314
rect 8496 734 8708 762
rect 10322 0 10378 800
<< via2 >>
rect 1991 10362 2047 10364
rect 2071 10362 2127 10364
rect 2151 10362 2207 10364
rect 2231 10362 2287 10364
rect 1991 10310 2037 10362
rect 2037 10310 2047 10362
rect 2071 10310 2101 10362
rect 2101 10310 2113 10362
rect 2113 10310 2127 10362
rect 2151 10310 2165 10362
rect 2165 10310 2177 10362
rect 2177 10310 2207 10362
rect 2231 10310 2241 10362
rect 2241 10310 2287 10362
rect 1991 10308 2047 10310
rect 2071 10308 2127 10310
rect 2151 10308 2207 10310
rect 2231 10308 2287 10310
rect 1398 10104 1454 10160
rect 2778 11872 2834 11928
rect 4061 10362 4117 10364
rect 4141 10362 4197 10364
rect 4221 10362 4277 10364
rect 4301 10362 4357 10364
rect 4061 10310 4107 10362
rect 4107 10310 4117 10362
rect 4141 10310 4171 10362
rect 4171 10310 4183 10362
rect 4183 10310 4197 10362
rect 4221 10310 4235 10362
rect 4235 10310 4247 10362
rect 4247 10310 4277 10362
rect 4301 10310 4311 10362
rect 4311 10310 4357 10362
rect 4061 10308 4117 10310
rect 4141 10308 4197 10310
rect 4221 10308 4277 10310
rect 4301 10308 4357 10310
rect 6131 10362 6187 10364
rect 6211 10362 6267 10364
rect 6291 10362 6347 10364
rect 6371 10362 6427 10364
rect 6131 10310 6177 10362
rect 6177 10310 6187 10362
rect 6211 10310 6241 10362
rect 6241 10310 6253 10362
rect 6253 10310 6267 10362
rect 6291 10310 6305 10362
rect 6305 10310 6317 10362
rect 6317 10310 6347 10362
rect 6371 10310 6381 10362
rect 6381 10310 6427 10362
rect 6131 10308 6187 10310
rect 6211 10308 6267 10310
rect 6291 10308 6347 10310
rect 6371 10308 6427 10310
rect 9310 11600 9366 11656
rect 8201 10362 8257 10364
rect 8281 10362 8337 10364
rect 8361 10362 8417 10364
rect 8441 10362 8497 10364
rect 8201 10310 8247 10362
rect 8247 10310 8257 10362
rect 8281 10310 8311 10362
rect 8311 10310 8323 10362
rect 8323 10310 8337 10362
rect 8361 10310 8375 10362
rect 8375 10310 8387 10362
rect 8387 10310 8417 10362
rect 8441 10310 8451 10362
rect 8451 10310 8497 10362
rect 8201 10308 8257 10310
rect 8281 10308 8337 10310
rect 8361 10308 8417 10310
rect 8441 10308 8497 10310
rect 938 8916 940 8936
rect 940 8916 992 8936
rect 992 8916 994 8936
rect 938 8880 994 8916
rect 1490 6840 1546 6896
rect 938 4800 994 4856
rect 938 3460 994 3496
rect 938 3440 940 3460
rect 940 3440 992 3460
rect 992 3440 994 3460
rect 1991 9274 2047 9276
rect 2071 9274 2127 9276
rect 2151 9274 2207 9276
rect 2231 9274 2287 9276
rect 1991 9222 2037 9274
rect 2037 9222 2047 9274
rect 2071 9222 2101 9274
rect 2101 9222 2113 9274
rect 2113 9222 2127 9274
rect 2151 9222 2165 9274
rect 2165 9222 2177 9274
rect 2177 9222 2207 9274
rect 2231 9222 2241 9274
rect 2241 9222 2287 9274
rect 1991 9220 2047 9222
rect 2071 9220 2127 9222
rect 2151 9220 2207 9222
rect 2231 9220 2287 9222
rect 1991 8186 2047 8188
rect 2071 8186 2127 8188
rect 2151 8186 2207 8188
rect 2231 8186 2287 8188
rect 1991 8134 2037 8186
rect 2037 8134 2047 8186
rect 2071 8134 2101 8186
rect 2101 8134 2113 8186
rect 2113 8134 2127 8186
rect 2151 8134 2165 8186
rect 2165 8134 2177 8186
rect 2177 8134 2207 8186
rect 2231 8134 2241 8186
rect 2241 8134 2287 8186
rect 1991 8132 2047 8134
rect 2071 8132 2127 8134
rect 2151 8132 2207 8134
rect 2231 8132 2287 8134
rect 1991 7098 2047 7100
rect 2071 7098 2127 7100
rect 2151 7098 2207 7100
rect 2231 7098 2287 7100
rect 1991 7046 2037 7098
rect 2037 7046 2047 7098
rect 2071 7046 2101 7098
rect 2101 7046 2113 7098
rect 2113 7046 2127 7098
rect 2151 7046 2165 7098
rect 2165 7046 2177 7098
rect 2177 7046 2207 7098
rect 2231 7046 2241 7098
rect 2241 7046 2287 7098
rect 1991 7044 2047 7046
rect 2071 7044 2127 7046
rect 2151 7044 2207 7046
rect 2231 7044 2287 7046
rect 1991 6010 2047 6012
rect 2071 6010 2127 6012
rect 2151 6010 2207 6012
rect 2231 6010 2287 6012
rect 1991 5958 2037 6010
rect 2037 5958 2047 6010
rect 2071 5958 2101 6010
rect 2101 5958 2113 6010
rect 2113 5958 2127 6010
rect 2151 5958 2165 6010
rect 2165 5958 2177 6010
rect 2177 5958 2207 6010
rect 2231 5958 2241 6010
rect 2241 5958 2287 6010
rect 1991 5956 2047 5958
rect 2071 5956 2127 5958
rect 2151 5956 2207 5958
rect 2231 5956 2287 5958
rect 1991 4922 2047 4924
rect 2071 4922 2127 4924
rect 2151 4922 2207 4924
rect 2231 4922 2287 4924
rect 1991 4870 2037 4922
rect 2037 4870 2047 4922
rect 2071 4870 2101 4922
rect 2101 4870 2113 4922
rect 2113 4870 2127 4922
rect 2151 4870 2165 4922
rect 2165 4870 2177 4922
rect 2177 4870 2207 4922
rect 2231 4870 2241 4922
rect 2241 4870 2287 4922
rect 1991 4868 2047 4870
rect 2071 4868 2127 4870
rect 2151 4868 2207 4870
rect 2231 4868 2287 4870
rect 1991 3834 2047 3836
rect 2071 3834 2127 3836
rect 2151 3834 2207 3836
rect 2231 3834 2287 3836
rect 1991 3782 2037 3834
rect 2037 3782 2047 3834
rect 2071 3782 2101 3834
rect 2101 3782 2113 3834
rect 2113 3782 2127 3834
rect 2151 3782 2165 3834
rect 2165 3782 2177 3834
rect 2177 3782 2207 3834
rect 2231 3782 2241 3834
rect 2241 3782 2287 3834
rect 1991 3780 2047 3782
rect 2071 3780 2127 3782
rect 2151 3780 2207 3782
rect 2231 3780 2287 3782
rect 2651 9818 2707 9820
rect 2731 9818 2787 9820
rect 2811 9818 2867 9820
rect 2891 9818 2947 9820
rect 2651 9766 2697 9818
rect 2697 9766 2707 9818
rect 2731 9766 2761 9818
rect 2761 9766 2773 9818
rect 2773 9766 2787 9818
rect 2811 9766 2825 9818
rect 2825 9766 2837 9818
rect 2837 9766 2867 9818
rect 2891 9766 2901 9818
rect 2901 9766 2947 9818
rect 2651 9764 2707 9766
rect 2731 9764 2787 9766
rect 2811 9764 2867 9766
rect 2891 9764 2947 9766
rect 3238 9580 3294 9616
rect 3238 9560 3240 9580
rect 3240 9560 3292 9580
rect 3292 9560 3294 9580
rect 2651 8730 2707 8732
rect 2731 8730 2787 8732
rect 2811 8730 2867 8732
rect 2891 8730 2947 8732
rect 2651 8678 2697 8730
rect 2697 8678 2707 8730
rect 2731 8678 2761 8730
rect 2761 8678 2773 8730
rect 2773 8678 2787 8730
rect 2811 8678 2825 8730
rect 2825 8678 2837 8730
rect 2837 8678 2867 8730
rect 2891 8678 2901 8730
rect 2901 8678 2947 8730
rect 2651 8676 2707 8678
rect 2731 8676 2787 8678
rect 2811 8676 2867 8678
rect 2891 8676 2947 8678
rect 2651 7642 2707 7644
rect 2731 7642 2787 7644
rect 2811 7642 2867 7644
rect 2891 7642 2947 7644
rect 2651 7590 2697 7642
rect 2697 7590 2707 7642
rect 2731 7590 2761 7642
rect 2761 7590 2773 7642
rect 2773 7590 2787 7642
rect 2811 7590 2825 7642
rect 2825 7590 2837 7642
rect 2837 7590 2867 7642
rect 2891 7590 2901 7642
rect 2901 7590 2947 7642
rect 2651 7588 2707 7590
rect 2731 7588 2787 7590
rect 2811 7588 2867 7590
rect 2891 7588 2947 7590
rect 2651 6554 2707 6556
rect 2731 6554 2787 6556
rect 2811 6554 2867 6556
rect 2891 6554 2947 6556
rect 2651 6502 2697 6554
rect 2697 6502 2707 6554
rect 2731 6502 2761 6554
rect 2761 6502 2773 6554
rect 2773 6502 2787 6554
rect 2811 6502 2825 6554
rect 2825 6502 2837 6554
rect 2837 6502 2867 6554
rect 2891 6502 2901 6554
rect 2901 6502 2947 6554
rect 2651 6500 2707 6502
rect 2731 6500 2787 6502
rect 2811 6500 2867 6502
rect 2891 6500 2947 6502
rect 2651 5466 2707 5468
rect 2731 5466 2787 5468
rect 2811 5466 2867 5468
rect 2891 5466 2947 5468
rect 2651 5414 2697 5466
rect 2697 5414 2707 5466
rect 2731 5414 2761 5466
rect 2761 5414 2773 5466
rect 2773 5414 2787 5466
rect 2811 5414 2825 5466
rect 2825 5414 2837 5466
rect 2837 5414 2867 5466
rect 2891 5414 2901 5466
rect 2901 5414 2947 5466
rect 2651 5412 2707 5414
rect 2731 5412 2787 5414
rect 2811 5412 2867 5414
rect 2891 5412 2947 5414
rect 4721 9818 4777 9820
rect 4801 9818 4857 9820
rect 4881 9818 4937 9820
rect 4961 9818 5017 9820
rect 4721 9766 4767 9818
rect 4767 9766 4777 9818
rect 4801 9766 4831 9818
rect 4831 9766 4843 9818
rect 4843 9766 4857 9818
rect 4881 9766 4895 9818
rect 4895 9766 4907 9818
rect 4907 9766 4937 9818
rect 4961 9766 4971 9818
rect 4971 9766 5017 9818
rect 4721 9764 4777 9766
rect 4801 9764 4857 9766
rect 4881 9764 4937 9766
rect 4961 9764 5017 9766
rect 4986 9580 5042 9616
rect 4986 9560 4988 9580
rect 4988 9560 5040 9580
rect 5040 9560 5042 9580
rect 4061 9274 4117 9276
rect 4141 9274 4197 9276
rect 4221 9274 4277 9276
rect 4301 9274 4357 9276
rect 4061 9222 4107 9274
rect 4107 9222 4117 9274
rect 4141 9222 4171 9274
rect 4171 9222 4183 9274
rect 4183 9222 4197 9274
rect 4221 9222 4235 9274
rect 4235 9222 4247 9274
rect 4247 9222 4277 9274
rect 4301 9222 4311 9274
rect 4311 9222 4357 9274
rect 4061 9220 4117 9222
rect 4141 9220 4197 9222
rect 4221 9220 4277 9222
rect 4301 9220 4357 9222
rect 5814 9560 5870 9616
rect 4061 8186 4117 8188
rect 4141 8186 4197 8188
rect 4221 8186 4277 8188
rect 4301 8186 4357 8188
rect 4061 8134 4107 8186
rect 4107 8134 4117 8186
rect 4141 8134 4171 8186
rect 4171 8134 4183 8186
rect 4183 8134 4197 8186
rect 4221 8134 4235 8186
rect 4235 8134 4247 8186
rect 4247 8134 4277 8186
rect 4301 8134 4311 8186
rect 4311 8134 4357 8186
rect 4061 8132 4117 8134
rect 4141 8132 4197 8134
rect 4221 8132 4277 8134
rect 4301 8132 4357 8134
rect 2651 4378 2707 4380
rect 2731 4378 2787 4380
rect 2811 4378 2867 4380
rect 2891 4378 2947 4380
rect 2651 4326 2697 4378
rect 2697 4326 2707 4378
rect 2731 4326 2761 4378
rect 2761 4326 2773 4378
rect 2773 4326 2787 4378
rect 2811 4326 2825 4378
rect 2825 4326 2837 4378
rect 2837 4326 2867 4378
rect 2891 4326 2901 4378
rect 2901 4326 2947 4378
rect 2651 4324 2707 4326
rect 2731 4324 2787 4326
rect 2811 4324 2867 4326
rect 2891 4324 2947 4326
rect 2651 3290 2707 3292
rect 2731 3290 2787 3292
rect 2811 3290 2867 3292
rect 2891 3290 2947 3292
rect 2651 3238 2697 3290
rect 2697 3238 2707 3290
rect 2731 3238 2761 3290
rect 2761 3238 2773 3290
rect 2773 3238 2787 3290
rect 2811 3238 2825 3290
rect 2825 3238 2837 3290
rect 2837 3238 2867 3290
rect 2891 3238 2901 3290
rect 2901 3238 2947 3290
rect 2651 3236 2707 3238
rect 2731 3236 2787 3238
rect 2811 3236 2867 3238
rect 2891 3236 2947 3238
rect 1991 2746 2047 2748
rect 2071 2746 2127 2748
rect 2151 2746 2207 2748
rect 2231 2746 2287 2748
rect 1991 2694 2037 2746
rect 2037 2694 2047 2746
rect 2071 2694 2101 2746
rect 2101 2694 2113 2746
rect 2113 2694 2127 2746
rect 2151 2694 2165 2746
rect 2165 2694 2177 2746
rect 2177 2694 2207 2746
rect 2231 2694 2241 2746
rect 2241 2694 2287 2746
rect 1991 2692 2047 2694
rect 2071 2692 2127 2694
rect 2151 2692 2207 2694
rect 2231 2692 2287 2694
rect 4061 7098 4117 7100
rect 4141 7098 4197 7100
rect 4221 7098 4277 7100
rect 4301 7098 4357 7100
rect 4061 7046 4107 7098
rect 4107 7046 4117 7098
rect 4141 7046 4171 7098
rect 4171 7046 4183 7098
rect 4183 7046 4197 7098
rect 4221 7046 4235 7098
rect 4235 7046 4247 7098
rect 4247 7046 4277 7098
rect 4301 7046 4311 7098
rect 4311 7046 4357 7098
rect 4061 7044 4117 7046
rect 4141 7044 4197 7046
rect 4221 7044 4277 7046
rect 4301 7044 4357 7046
rect 4721 8730 4777 8732
rect 4801 8730 4857 8732
rect 4881 8730 4937 8732
rect 4961 8730 5017 8732
rect 4721 8678 4767 8730
rect 4767 8678 4777 8730
rect 4801 8678 4831 8730
rect 4831 8678 4843 8730
rect 4843 8678 4857 8730
rect 4881 8678 4895 8730
rect 4895 8678 4907 8730
rect 4907 8678 4937 8730
rect 4961 8678 4971 8730
rect 4971 8678 5017 8730
rect 4721 8676 4777 8678
rect 4801 8676 4857 8678
rect 4881 8676 4937 8678
rect 4961 8676 5017 8678
rect 4721 7642 4777 7644
rect 4801 7642 4857 7644
rect 4881 7642 4937 7644
rect 4961 7642 5017 7644
rect 4721 7590 4767 7642
rect 4767 7590 4777 7642
rect 4801 7590 4831 7642
rect 4831 7590 4843 7642
rect 4843 7590 4857 7642
rect 4881 7590 4895 7642
rect 4895 7590 4907 7642
rect 4907 7590 4937 7642
rect 4961 7590 4971 7642
rect 4971 7590 5017 7642
rect 4721 7588 4777 7590
rect 4801 7588 4857 7590
rect 4881 7588 4937 7590
rect 4961 7588 5017 7590
rect 4061 6010 4117 6012
rect 4141 6010 4197 6012
rect 4221 6010 4277 6012
rect 4301 6010 4357 6012
rect 4061 5958 4107 6010
rect 4107 5958 4117 6010
rect 4141 5958 4171 6010
rect 4171 5958 4183 6010
rect 4183 5958 4197 6010
rect 4221 5958 4235 6010
rect 4235 5958 4247 6010
rect 4247 5958 4277 6010
rect 4301 5958 4311 6010
rect 4311 5958 4357 6010
rect 4061 5956 4117 5958
rect 4141 5956 4197 5958
rect 4221 5956 4277 5958
rect 4301 5956 4357 5958
rect 4061 4922 4117 4924
rect 4141 4922 4197 4924
rect 4221 4922 4277 4924
rect 4301 4922 4357 4924
rect 4061 4870 4107 4922
rect 4107 4870 4117 4922
rect 4141 4870 4171 4922
rect 4171 4870 4183 4922
rect 4183 4870 4197 4922
rect 4221 4870 4235 4922
rect 4235 4870 4247 4922
rect 4247 4870 4277 4922
rect 4301 4870 4311 4922
rect 4311 4870 4357 4922
rect 4061 4868 4117 4870
rect 4141 4868 4197 4870
rect 4221 4868 4277 4870
rect 4301 4868 4357 4870
rect 4061 3834 4117 3836
rect 4141 3834 4197 3836
rect 4221 3834 4277 3836
rect 4301 3834 4357 3836
rect 4061 3782 4107 3834
rect 4107 3782 4117 3834
rect 4141 3782 4171 3834
rect 4171 3782 4183 3834
rect 4183 3782 4197 3834
rect 4221 3782 4235 3834
rect 4235 3782 4247 3834
rect 4247 3782 4277 3834
rect 4301 3782 4311 3834
rect 4311 3782 4357 3834
rect 4061 3780 4117 3782
rect 4141 3780 4197 3782
rect 4221 3780 4277 3782
rect 4301 3780 4357 3782
rect 4721 6554 4777 6556
rect 4801 6554 4857 6556
rect 4881 6554 4937 6556
rect 4961 6554 5017 6556
rect 4721 6502 4767 6554
rect 4767 6502 4777 6554
rect 4801 6502 4831 6554
rect 4831 6502 4843 6554
rect 4843 6502 4857 6554
rect 4881 6502 4895 6554
rect 4895 6502 4907 6554
rect 4907 6502 4937 6554
rect 4961 6502 4971 6554
rect 4971 6502 5017 6554
rect 4721 6500 4777 6502
rect 4801 6500 4857 6502
rect 4881 6500 4937 6502
rect 4961 6500 5017 6502
rect 4721 5466 4777 5468
rect 4801 5466 4857 5468
rect 4881 5466 4937 5468
rect 4961 5466 5017 5468
rect 4721 5414 4767 5466
rect 4767 5414 4777 5466
rect 4801 5414 4831 5466
rect 4831 5414 4843 5466
rect 4843 5414 4857 5466
rect 4881 5414 4895 5466
rect 4895 5414 4907 5466
rect 4907 5414 4937 5466
rect 4961 5414 4971 5466
rect 4971 5414 5017 5466
rect 4721 5412 4777 5414
rect 4801 5412 4857 5414
rect 4881 5412 4937 5414
rect 4961 5412 5017 5414
rect 6131 9274 6187 9276
rect 6211 9274 6267 9276
rect 6291 9274 6347 9276
rect 6371 9274 6427 9276
rect 6131 9222 6177 9274
rect 6177 9222 6187 9274
rect 6211 9222 6241 9274
rect 6241 9222 6253 9274
rect 6253 9222 6267 9274
rect 6291 9222 6305 9274
rect 6305 9222 6317 9274
rect 6317 9222 6347 9274
rect 6371 9222 6381 9274
rect 6381 9222 6427 9274
rect 6131 9220 6187 9222
rect 6211 9220 6267 9222
rect 6291 9220 6347 9222
rect 6371 9220 6427 9222
rect 6131 8186 6187 8188
rect 6211 8186 6267 8188
rect 6291 8186 6347 8188
rect 6371 8186 6427 8188
rect 6131 8134 6177 8186
rect 6177 8134 6187 8186
rect 6211 8134 6241 8186
rect 6241 8134 6253 8186
rect 6253 8134 6267 8186
rect 6291 8134 6305 8186
rect 6305 8134 6317 8186
rect 6317 8134 6347 8186
rect 6371 8134 6381 8186
rect 6381 8134 6427 8186
rect 6131 8132 6187 8134
rect 6211 8132 6267 8134
rect 6291 8132 6347 8134
rect 6371 8132 6427 8134
rect 4721 4378 4777 4380
rect 4801 4378 4857 4380
rect 4881 4378 4937 4380
rect 4961 4378 5017 4380
rect 4721 4326 4767 4378
rect 4767 4326 4777 4378
rect 4801 4326 4831 4378
rect 4831 4326 4843 4378
rect 4843 4326 4857 4378
rect 4881 4326 4895 4378
rect 4895 4326 4907 4378
rect 4907 4326 4937 4378
rect 4961 4326 4971 4378
rect 4971 4326 5017 4378
rect 4721 4324 4777 4326
rect 4801 4324 4857 4326
rect 4881 4324 4937 4326
rect 4961 4324 5017 4326
rect 4721 3290 4777 3292
rect 4801 3290 4857 3292
rect 4881 3290 4937 3292
rect 4961 3290 5017 3292
rect 4721 3238 4767 3290
rect 4767 3238 4777 3290
rect 4801 3238 4831 3290
rect 4831 3238 4843 3290
rect 4843 3238 4857 3290
rect 4881 3238 4895 3290
rect 4895 3238 4907 3290
rect 4907 3238 4937 3290
rect 4961 3238 4971 3290
rect 4971 3238 5017 3290
rect 4721 3236 4777 3238
rect 4801 3236 4857 3238
rect 4881 3236 4937 3238
rect 4961 3236 5017 3238
rect 4061 2746 4117 2748
rect 4141 2746 4197 2748
rect 4221 2746 4277 2748
rect 4301 2746 4357 2748
rect 4061 2694 4107 2746
rect 4107 2694 4117 2746
rect 4141 2694 4171 2746
rect 4171 2694 4183 2746
rect 4183 2694 4197 2746
rect 4221 2694 4235 2746
rect 4235 2694 4247 2746
rect 4247 2694 4277 2746
rect 4301 2694 4311 2746
rect 4311 2694 4357 2746
rect 4061 2692 4117 2694
rect 4141 2692 4197 2694
rect 4221 2692 4277 2694
rect 4301 2692 4357 2694
rect 1214 1400 1270 1456
rect 6131 7098 6187 7100
rect 6211 7098 6267 7100
rect 6291 7098 6347 7100
rect 6371 7098 6427 7100
rect 6131 7046 6177 7098
rect 6177 7046 6187 7098
rect 6211 7046 6241 7098
rect 6241 7046 6253 7098
rect 6253 7046 6267 7098
rect 6291 7046 6305 7098
rect 6305 7046 6317 7098
rect 6317 7046 6347 7098
rect 6371 7046 6381 7098
rect 6381 7046 6427 7098
rect 6131 7044 6187 7046
rect 6211 7044 6267 7046
rect 6291 7044 6347 7046
rect 6371 7044 6427 7046
rect 6791 9818 6847 9820
rect 6871 9818 6927 9820
rect 6951 9818 7007 9820
rect 7031 9818 7087 9820
rect 6791 9766 6837 9818
rect 6837 9766 6847 9818
rect 6871 9766 6901 9818
rect 6901 9766 6913 9818
rect 6913 9766 6927 9818
rect 6951 9766 6965 9818
rect 6965 9766 6977 9818
rect 6977 9766 7007 9818
rect 7031 9766 7041 9818
rect 7041 9766 7087 9818
rect 6791 9764 6847 9766
rect 6871 9764 6927 9766
rect 6951 9764 7007 9766
rect 7031 9764 7087 9766
rect 6791 8730 6847 8732
rect 6871 8730 6927 8732
rect 6951 8730 7007 8732
rect 7031 8730 7087 8732
rect 6791 8678 6837 8730
rect 6837 8678 6847 8730
rect 6871 8678 6901 8730
rect 6901 8678 6913 8730
rect 6913 8678 6927 8730
rect 6951 8678 6965 8730
rect 6965 8678 6977 8730
rect 6977 8678 7007 8730
rect 7031 8678 7041 8730
rect 7041 8678 7087 8730
rect 6791 8676 6847 8678
rect 6871 8676 6927 8678
rect 6951 8676 7007 8678
rect 7031 8676 7087 8678
rect 6791 7642 6847 7644
rect 6871 7642 6927 7644
rect 6951 7642 7007 7644
rect 7031 7642 7087 7644
rect 6791 7590 6837 7642
rect 6837 7590 6847 7642
rect 6871 7590 6901 7642
rect 6901 7590 6913 7642
rect 6913 7590 6927 7642
rect 6951 7590 6965 7642
rect 6965 7590 6977 7642
rect 6977 7590 7007 7642
rect 7031 7590 7041 7642
rect 7041 7590 7087 7642
rect 6791 7588 6847 7590
rect 6871 7588 6927 7590
rect 6951 7588 7007 7590
rect 7031 7588 7087 7590
rect 6791 6554 6847 6556
rect 6871 6554 6927 6556
rect 6951 6554 7007 6556
rect 7031 6554 7087 6556
rect 6791 6502 6837 6554
rect 6837 6502 6847 6554
rect 6871 6502 6901 6554
rect 6901 6502 6913 6554
rect 6913 6502 6927 6554
rect 6951 6502 6965 6554
rect 6965 6502 6977 6554
rect 6977 6502 7007 6554
rect 7031 6502 7041 6554
rect 7041 6502 7087 6554
rect 6791 6500 6847 6502
rect 6871 6500 6927 6502
rect 6951 6500 7007 6502
rect 7031 6500 7087 6502
rect 6131 6010 6187 6012
rect 6211 6010 6267 6012
rect 6291 6010 6347 6012
rect 6371 6010 6427 6012
rect 6131 5958 6177 6010
rect 6177 5958 6187 6010
rect 6211 5958 6241 6010
rect 6241 5958 6253 6010
rect 6253 5958 6267 6010
rect 6291 5958 6305 6010
rect 6305 5958 6317 6010
rect 6317 5958 6347 6010
rect 6371 5958 6381 6010
rect 6381 5958 6427 6010
rect 6131 5956 6187 5958
rect 6211 5956 6267 5958
rect 6291 5956 6347 5958
rect 6371 5956 6427 5958
rect 6131 4922 6187 4924
rect 6211 4922 6267 4924
rect 6291 4922 6347 4924
rect 6371 4922 6427 4924
rect 6131 4870 6177 4922
rect 6177 4870 6187 4922
rect 6211 4870 6241 4922
rect 6241 4870 6253 4922
rect 6253 4870 6267 4922
rect 6291 4870 6305 4922
rect 6305 4870 6317 4922
rect 6317 4870 6347 4922
rect 6371 4870 6381 4922
rect 6381 4870 6427 4922
rect 6131 4868 6187 4870
rect 6211 4868 6267 4870
rect 6291 4868 6347 4870
rect 6371 4868 6427 4870
rect 6131 3834 6187 3836
rect 6211 3834 6267 3836
rect 6291 3834 6347 3836
rect 6371 3834 6427 3836
rect 6131 3782 6177 3834
rect 6177 3782 6187 3834
rect 6211 3782 6241 3834
rect 6241 3782 6253 3834
rect 6253 3782 6267 3834
rect 6291 3782 6305 3834
rect 6305 3782 6317 3834
rect 6317 3782 6347 3834
rect 6371 3782 6381 3834
rect 6381 3782 6427 3834
rect 6131 3780 6187 3782
rect 6211 3780 6267 3782
rect 6291 3780 6347 3782
rect 6371 3780 6427 3782
rect 6791 5466 6847 5468
rect 6871 5466 6927 5468
rect 6951 5466 7007 5468
rect 7031 5466 7087 5468
rect 6791 5414 6837 5466
rect 6837 5414 6847 5466
rect 6871 5414 6901 5466
rect 6901 5414 6913 5466
rect 6913 5414 6927 5466
rect 6951 5414 6965 5466
rect 6965 5414 6977 5466
rect 6977 5414 7007 5466
rect 7031 5414 7041 5466
rect 7041 5414 7087 5466
rect 6791 5412 6847 5414
rect 6871 5412 6927 5414
rect 6951 5412 7007 5414
rect 7031 5412 7087 5414
rect 7378 9580 7434 9616
rect 7378 9560 7380 9580
rect 7380 9560 7432 9580
rect 7432 9560 7434 9580
rect 6131 2746 6187 2748
rect 6211 2746 6267 2748
rect 6291 2746 6347 2748
rect 6371 2746 6427 2748
rect 6131 2694 6177 2746
rect 6177 2694 6187 2746
rect 6211 2694 6241 2746
rect 6241 2694 6253 2746
rect 6253 2694 6267 2746
rect 6291 2694 6305 2746
rect 6305 2694 6317 2746
rect 6317 2694 6347 2746
rect 6371 2694 6381 2746
rect 6381 2694 6427 2746
rect 6131 2692 6187 2694
rect 6211 2692 6267 2694
rect 6291 2692 6347 2694
rect 6371 2692 6427 2694
rect 6791 4378 6847 4380
rect 6871 4378 6927 4380
rect 6951 4378 7007 4380
rect 7031 4378 7087 4380
rect 6791 4326 6837 4378
rect 6837 4326 6847 4378
rect 6871 4326 6901 4378
rect 6901 4326 6913 4378
rect 6913 4326 6927 4378
rect 6951 4326 6965 4378
rect 6965 4326 6977 4378
rect 6977 4326 7007 4378
rect 7031 4326 7041 4378
rect 7041 4326 7087 4378
rect 6791 4324 6847 4326
rect 6871 4324 6927 4326
rect 6951 4324 7007 4326
rect 7031 4324 7087 4326
rect 6791 3290 6847 3292
rect 6871 3290 6927 3292
rect 6951 3290 7007 3292
rect 7031 3290 7087 3292
rect 6791 3238 6837 3290
rect 6837 3238 6847 3290
rect 6871 3238 6901 3290
rect 6901 3238 6913 3290
rect 6913 3238 6927 3290
rect 6951 3238 6965 3290
rect 6965 3238 6977 3290
rect 6977 3238 7007 3290
rect 7031 3238 7041 3290
rect 7041 3238 7087 3290
rect 6791 3236 6847 3238
rect 6871 3236 6927 3238
rect 6951 3236 7007 3238
rect 7031 3236 7087 3238
rect 8201 9274 8257 9276
rect 8281 9274 8337 9276
rect 8361 9274 8417 9276
rect 8441 9274 8497 9276
rect 8201 9222 8247 9274
rect 8247 9222 8257 9274
rect 8281 9222 8311 9274
rect 8311 9222 8323 9274
rect 8323 9222 8337 9274
rect 8361 9222 8375 9274
rect 8375 9222 8387 9274
rect 8387 9222 8417 9274
rect 8441 9222 8451 9274
rect 8451 9222 8497 9274
rect 8201 9220 8257 9222
rect 8281 9220 8337 9222
rect 8361 9220 8417 9222
rect 8441 9220 8497 9222
rect 8861 9818 8917 9820
rect 8941 9818 8997 9820
rect 9021 9818 9077 9820
rect 9101 9818 9157 9820
rect 8861 9766 8907 9818
rect 8907 9766 8917 9818
rect 8941 9766 8971 9818
rect 8971 9766 8983 9818
rect 8983 9766 8997 9818
rect 9021 9766 9035 9818
rect 9035 9766 9047 9818
rect 9047 9766 9077 9818
rect 9101 9766 9111 9818
rect 9111 9766 9157 9818
rect 8861 9764 8917 9766
rect 8941 9764 8997 9766
rect 9021 9764 9077 9766
rect 9101 9764 9157 9766
rect 9402 10240 9458 10296
rect 8861 8730 8917 8732
rect 8941 8730 8997 8732
rect 9021 8730 9077 8732
rect 9101 8730 9157 8732
rect 8861 8678 8907 8730
rect 8907 8678 8917 8730
rect 8941 8678 8971 8730
rect 8971 8678 8983 8730
rect 8983 8678 8997 8730
rect 9021 8678 9035 8730
rect 9035 8678 9047 8730
rect 9047 8678 9077 8730
rect 9101 8678 9111 8730
rect 9111 8678 9157 8730
rect 8861 8676 8917 8678
rect 8941 8676 8997 8678
rect 9021 8676 9077 8678
rect 9101 8676 9157 8678
rect 8201 8186 8257 8188
rect 8281 8186 8337 8188
rect 8361 8186 8417 8188
rect 8441 8186 8497 8188
rect 8201 8134 8247 8186
rect 8247 8134 8257 8186
rect 8281 8134 8311 8186
rect 8311 8134 8323 8186
rect 8323 8134 8337 8186
rect 8361 8134 8375 8186
rect 8375 8134 8387 8186
rect 8387 8134 8417 8186
rect 8441 8134 8451 8186
rect 8451 8134 8497 8186
rect 8201 8132 8257 8134
rect 8281 8132 8337 8134
rect 8361 8132 8417 8134
rect 8441 8132 8497 8134
rect 9034 8200 9090 8256
rect 8861 7642 8917 7644
rect 8941 7642 8997 7644
rect 9021 7642 9077 7644
rect 9101 7642 9157 7644
rect 8861 7590 8907 7642
rect 8907 7590 8917 7642
rect 8941 7590 8971 7642
rect 8971 7590 8983 7642
rect 8983 7590 8997 7642
rect 9021 7590 9035 7642
rect 9035 7590 9047 7642
rect 9047 7590 9077 7642
rect 9101 7590 9111 7642
rect 9111 7590 9157 7642
rect 8861 7588 8917 7590
rect 8941 7588 8997 7590
rect 9021 7588 9077 7590
rect 9101 7588 9157 7590
rect 8201 7098 8257 7100
rect 8281 7098 8337 7100
rect 8361 7098 8417 7100
rect 8441 7098 8497 7100
rect 8201 7046 8247 7098
rect 8247 7046 8257 7098
rect 8281 7046 8311 7098
rect 8311 7046 8323 7098
rect 8323 7046 8337 7098
rect 8361 7046 8375 7098
rect 8375 7046 8387 7098
rect 8387 7046 8417 7098
rect 8441 7046 8451 7098
rect 8451 7046 8497 7098
rect 8201 7044 8257 7046
rect 8281 7044 8337 7046
rect 8361 7044 8417 7046
rect 8441 7044 8497 7046
rect 8861 6554 8917 6556
rect 8941 6554 8997 6556
rect 9021 6554 9077 6556
rect 9101 6554 9157 6556
rect 8861 6502 8907 6554
rect 8907 6502 8917 6554
rect 8941 6502 8971 6554
rect 8971 6502 8983 6554
rect 8983 6502 8997 6554
rect 9021 6502 9035 6554
rect 9035 6502 9047 6554
rect 9047 6502 9077 6554
rect 9101 6502 9111 6554
rect 9111 6502 9157 6554
rect 8861 6500 8917 6502
rect 8941 6500 8997 6502
rect 9021 6500 9077 6502
rect 9101 6500 9157 6502
rect 8201 6010 8257 6012
rect 8281 6010 8337 6012
rect 8361 6010 8417 6012
rect 8441 6010 8497 6012
rect 8201 5958 8247 6010
rect 8247 5958 8257 6010
rect 8281 5958 8311 6010
rect 8311 5958 8323 6010
rect 8323 5958 8337 6010
rect 8361 5958 8375 6010
rect 8375 5958 8387 6010
rect 8387 5958 8417 6010
rect 8441 5958 8451 6010
rect 8451 5958 8497 6010
rect 8201 5956 8257 5958
rect 8281 5956 8337 5958
rect 8361 5956 8417 5958
rect 8441 5956 8497 5958
rect 8201 4922 8257 4924
rect 8281 4922 8337 4924
rect 8361 4922 8417 4924
rect 8441 4922 8497 4924
rect 8201 4870 8247 4922
rect 8247 4870 8257 4922
rect 8281 4870 8311 4922
rect 8311 4870 8323 4922
rect 8323 4870 8337 4922
rect 8361 4870 8375 4922
rect 8375 4870 8387 4922
rect 8387 4870 8417 4922
rect 8441 4870 8451 4922
rect 8451 4870 8497 4922
rect 8201 4868 8257 4870
rect 8281 4868 8337 4870
rect 8361 4868 8417 4870
rect 8441 4868 8497 4870
rect 8201 3834 8257 3836
rect 8281 3834 8337 3836
rect 8361 3834 8417 3836
rect 8441 3834 8497 3836
rect 8201 3782 8247 3834
rect 8247 3782 8257 3834
rect 8281 3782 8311 3834
rect 8311 3782 8323 3834
rect 8323 3782 8337 3834
rect 8361 3782 8375 3834
rect 8375 3782 8387 3834
rect 8387 3782 8417 3834
rect 8441 3782 8451 3834
rect 8451 3782 8497 3834
rect 8201 3780 8257 3782
rect 8281 3780 8337 3782
rect 8361 3780 8417 3782
rect 8441 3780 8497 3782
rect 8666 6160 8722 6216
rect 8861 5466 8917 5468
rect 8941 5466 8997 5468
rect 9021 5466 9077 5468
rect 9101 5466 9157 5468
rect 8861 5414 8907 5466
rect 8907 5414 8917 5466
rect 8941 5414 8971 5466
rect 8971 5414 8983 5466
rect 8983 5414 8997 5466
rect 9021 5414 9035 5466
rect 9035 5414 9047 5466
rect 9047 5414 9077 5466
rect 9101 5414 9111 5466
rect 9111 5414 9157 5466
rect 8861 5412 8917 5414
rect 8941 5412 8997 5414
rect 9021 5412 9077 5414
rect 9101 5412 9157 5414
rect 9034 4800 9090 4856
rect 8861 4378 8917 4380
rect 8941 4378 8997 4380
rect 9021 4378 9077 4380
rect 9101 4378 9157 4380
rect 8861 4326 8907 4378
rect 8907 4326 8917 4378
rect 8941 4326 8971 4378
rect 8971 4326 8983 4378
rect 8983 4326 8997 4378
rect 9021 4326 9035 4378
rect 9035 4326 9047 4378
rect 9047 4326 9077 4378
rect 9101 4326 9111 4378
rect 9111 4326 9157 4378
rect 8861 4324 8917 4326
rect 8941 4324 8997 4326
rect 9021 4324 9077 4326
rect 9101 4324 9157 4326
rect 2651 2202 2707 2204
rect 2731 2202 2787 2204
rect 2811 2202 2867 2204
rect 2891 2202 2947 2204
rect 2651 2150 2697 2202
rect 2697 2150 2707 2202
rect 2731 2150 2761 2202
rect 2761 2150 2773 2202
rect 2773 2150 2787 2202
rect 2811 2150 2825 2202
rect 2825 2150 2837 2202
rect 2837 2150 2867 2202
rect 2891 2150 2901 2202
rect 2901 2150 2947 2202
rect 2651 2148 2707 2150
rect 2731 2148 2787 2150
rect 2811 2148 2867 2150
rect 2891 2148 2947 2150
rect 4721 2202 4777 2204
rect 4801 2202 4857 2204
rect 4881 2202 4937 2204
rect 4961 2202 5017 2204
rect 4721 2150 4767 2202
rect 4767 2150 4777 2202
rect 4801 2150 4831 2202
rect 4831 2150 4843 2202
rect 4843 2150 4857 2202
rect 4881 2150 4895 2202
rect 4895 2150 4907 2202
rect 4907 2150 4937 2202
rect 4961 2150 4971 2202
rect 4971 2150 5017 2202
rect 4721 2148 4777 2150
rect 4801 2148 4857 2150
rect 4881 2148 4937 2150
rect 4961 2148 5017 2150
rect 6791 2202 6847 2204
rect 6871 2202 6927 2204
rect 6951 2202 7007 2204
rect 7031 2202 7087 2204
rect 6791 2150 6837 2202
rect 6837 2150 6847 2202
rect 6871 2150 6901 2202
rect 6901 2150 6913 2202
rect 6913 2150 6927 2202
rect 6951 2150 6965 2202
rect 6965 2150 6977 2202
rect 6977 2150 7007 2202
rect 7031 2150 7041 2202
rect 7041 2150 7087 2202
rect 6791 2148 6847 2150
rect 6871 2148 6927 2150
rect 6951 2148 7007 2150
rect 7031 2148 7087 2150
rect 8201 2746 8257 2748
rect 8281 2746 8337 2748
rect 8361 2746 8417 2748
rect 8441 2746 8497 2748
rect 8201 2694 8247 2746
rect 8247 2694 8257 2746
rect 8281 2694 8311 2746
rect 8311 2694 8323 2746
rect 8323 2694 8337 2746
rect 8361 2694 8375 2746
rect 8375 2694 8387 2746
rect 8387 2694 8417 2746
rect 8441 2694 8451 2746
rect 8451 2694 8497 2746
rect 8201 2692 8257 2694
rect 8281 2692 8337 2694
rect 8361 2692 8417 2694
rect 8441 2692 8497 2694
rect 8022 720 8078 776
rect 8861 3290 8917 3292
rect 8941 3290 8997 3292
rect 9021 3290 9077 3292
rect 9101 3290 9157 3292
rect 8861 3238 8907 3290
rect 8907 3238 8917 3290
rect 8941 3238 8971 3290
rect 8971 3238 8983 3290
rect 8983 3238 8997 3290
rect 9021 3238 9035 3290
rect 9035 3238 9047 3290
rect 9047 3238 9077 3290
rect 9101 3238 9111 3290
rect 9111 3238 9157 3290
rect 8861 3236 8917 3238
rect 8941 3236 8997 3238
rect 9021 3236 9077 3238
rect 9101 3236 9157 3238
rect 9402 2760 9458 2816
rect 8861 2202 8917 2204
rect 8941 2202 8997 2204
rect 9021 2202 9077 2204
rect 9101 2202 9157 2204
rect 8861 2150 8907 2202
rect 8907 2150 8917 2202
rect 8941 2150 8971 2202
rect 8971 2150 8983 2202
rect 8983 2150 8997 2202
rect 9021 2150 9035 2202
rect 9035 2150 9047 2202
rect 9047 2150 9077 2202
rect 9101 2150 9111 2202
rect 9111 2150 9157 2202
rect 8861 2148 8917 2150
rect 8941 2148 8997 2150
rect 9021 2148 9077 2150
rect 9101 2148 9157 2150
<< metal3 >>
rect 0 12338 800 12368
rect 0 12278 1226 12338
rect 0 12248 800 12278
rect 1166 11930 1226 12278
rect 2773 11930 2839 11933
rect 1166 11928 2839 11930
rect 1166 11872 2778 11928
rect 2834 11872 2839 11928
rect 1166 11870 2839 11872
rect 2773 11867 2839 11870
rect 9305 11658 9371 11661
rect 9767 11658 10567 11688
rect 9305 11656 10567 11658
rect 9305 11600 9310 11656
rect 9366 11600 10567 11656
rect 9305 11598 10567 11600
rect 9305 11595 9371 11598
rect 9767 11568 10567 11598
rect 1981 10368 2297 10369
rect 0 10298 800 10328
rect 1981 10304 1987 10368
rect 2051 10304 2067 10368
rect 2131 10304 2147 10368
rect 2211 10304 2227 10368
rect 2291 10304 2297 10368
rect 1981 10303 2297 10304
rect 4051 10368 4367 10369
rect 4051 10304 4057 10368
rect 4121 10304 4137 10368
rect 4201 10304 4217 10368
rect 4281 10304 4297 10368
rect 4361 10304 4367 10368
rect 4051 10303 4367 10304
rect 6121 10368 6437 10369
rect 6121 10304 6127 10368
rect 6191 10304 6207 10368
rect 6271 10304 6287 10368
rect 6351 10304 6367 10368
rect 6431 10304 6437 10368
rect 6121 10303 6437 10304
rect 8191 10368 8507 10369
rect 8191 10304 8197 10368
rect 8261 10304 8277 10368
rect 8341 10304 8357 10368
rect 8421 10304 8437 10368
rect 8501 10304 8507 10368
rect 8191 10303 8507 10304
rect 9397 10298 9463 10301
rect 9767 10298 10567 10328
rect 0 10238 1594 10298
rect 0 10208 800 10238
rect 1393 10162 1459 10165
rect 1534 10162 1594 10238
rect 9397 10296 10567 10298
rect 9397 10240 9402 10296
rect 9458 10240 10567 10296
rect 9397 10238 10567 10240
rect 9397 10235 9463 10238
rect 9767 10208 10567 10238
rect 1393 10160 1594 10162
rect 1393 10104 1398 10160
rect 1454 10104 1594 10160
rect 1393 10102 1594 10104
rect 1393 10099 1459 10102
rect 2641 9824 2957 9825
rect 2641 9760 2647 9824
rect 2711 9760 2727 9824
rect 2791 9760 2807 9824
rect 2871 9760 2887 9824
rect 2951 9760 2957 9824
rect 2641 9759 2957 9760
rect 4711 9824 5027 9825
rect 4711 9760 4717 9824
rect 4781 9760 4797 9824
rect 4861 9760 4877 9824
rect 4941 9760 4957 9824
rect 5021 9760 5027 9824
rect 4711 9759 5027 9760
rect 6781 9824 7097 9825
rect 6781 9760 6787 9824
rect 6851 9760 6867 9824
rect 6931 9760 6947 9824
rect 7011 9760 7027 9824
rect 7091 9760 7097 9824
rect 6781 9759 7097 9760
rect 8851 9824 9167 9825
rect 8851 9760 8857 9824
rect 8921 9760 8937 9824
rect 9001 9760 9017 9824
rect 9081 9760 9097 9824
rect 9161 9760 9167 9824
rect 8851 9759 9167 9760
rect 3233 9618 3299 9621
rect 4981 9618 5047 9621
rect 3233 9616 5047 9618
rect 3233 9560 3238 9616
rect 3294 9560 4986 9616
rect 5042 9560 5047 9616
rect 3233 9558 5047 9560
rect 3233 9555 3299 9558
rect 4981 9555 5047 9558
rect 5809 9618 5875 9621
rect 7373 9618 7439 9621
rect 5809 9616 7439 9618
rect 5809 9560 5814 9616
rect 5870 9560 7378 9616
rect 7434 9560 7439 9616
rect 5809 9558 7439 9560
rect 5809 9555 5875 9558
rect 7373 9555 7439 9558
rect 1981 9280 2297 9281
rect 1981 9216 1987 9280
rect 2051 9216 2067 9280
rect 2131 9216 2147 9280
rect 2211 9216 2227 9280
rect 2291 9216 2297 9280
rect 1981 9215 2297 9216
rect 4051 9280 4367 9281
rect 4051 9216 4057 9280
rect 4121 9216 4137 9280
rect 4201 9216 4217 9280
rect 4281 9216 4297 9280
rect 4361 9216 4367 9280
rect 4051 9215 4367 9216
rect 6121 9280 6437 9281
rect 6121 9216 6127 9280
rect 6191 9216 6207 9280
rect 6271 9216 6287 9280
rect 6351 9216 6367 9280
rect 6431 9216 6437 9280
rect 6121 9215 6437 9216
rect 8191 9280 8507 9281
rect 8191 9216 8197 9280
rect 8261 9216 8277 9280
rect 8341 9216 8357 9280
rect 8421 9216 8437 9280
rect 8501 9216 8507 9280
rect 8191 9215 8507 9216
rect 0 8938 800 8968
rect 933 8938 999 8941
rect 0 8936 999 8938
rect 0 8880 938 8936
rect 994 8880 999 8936
rect 0 8878 999 8880
rect 0 8848 800 8878
rect 933 8875 999 8878
rect 2641 8736 2957 8737
rect 2641 8672 2647 8736
rect 2711 8672 2727 8736
rect 2791 8672 2807 8736
rect 2871 8672 2887 8736
rect 2951 8672 2957 8736
rect 2641 8671 2957 8672
rect 4711 8736 5027 8737
rect 4711 8672 4717 8736
rect 4781 8672 4797 8736
rect 4861 8672 4877 8736
rect 4941 8672 4957 8736
rect 5021 8672 5027 8736
rect 4711 8671 5027 8672
rect 6781 8736 7097 8737
rect 6781 8672 6787 8736
rect 6851 8672 6867 8736
rect 6931 8672 6947 8736
rect 7011 8672 7027 8736
rect 7091 8672 7097 8736
rect 6781 8671 7097 8672
rect 8851 8736 9167 8737
rect 8851 8672 8857 8736
rect 8921 8672 8937 8736
rect 9001 8672 9017 8736
rect 9081 8672 9097 8736
rect 9161 8672 9167 8736
rect 8851 8671 9167 8672
rect 9029 8258 9095 8261
rect 9767 8258 10567 8288
rect 9029 8256 10567 8258
rect 9029 8200 9034 8256
rect 9090 8200 10567 8256
rect 9029 8198 10567 8200
rect 9029 8195 9095 8198
rect 1981 8192 2297 8193
rect 1981 8128 1987 8192
rect 2051 8128 2067 8192
rect 2131 8128 2147 8192
rect 2211 8128 2227 8192
rect 2291 8128 2297 8192
rect 1981 8127 2297 8128
rect 4051 8192 4367 8193
rect 4051 8128 4057 8192
rect 4121 8128 4137 8192
rect 4201 8128 4217 8192
rect 4281 8128 4297 8192
rect 4361 8128 4367 8192
rect 4051 8127 4367 8128
rect 6121 8192 6437 8193
rect 6121 8128 6127 8192
rect 6191 8128 6207 8192
rect 6271 8128 6287 8192
rect 6351 8128 6367 8192
rect 6431 8128 6437 8192
rect 6121 8127 6437 8128
rect 8191 8192 8507 8193
rect 8191 8128 8197 8192
rect 8261 8128 8277 8192
rect 8341 8128 8357 8192
rect 8421 8128 8437 8192
rect 8501 8128 8507 8192
rect 9767 8168 10567 8198
rect 8191 8127 8507 8128
rect 2641 7648 2957 7649
rect 2641 7584 2647 7648
rect 2711 7584 2727 7648
rect 2791 7584 2807 7648
rect 2871 7584 2887 7648
rect 2951 7584 2957 7648
rect 2641 7583 2957 7584
rect 4711 7648 5027 7649
rect 4711 7584 4717 7648
rect 4781 7584 4797 7648
rect 4861 7584 4877 7648
rect 4941 7584 4957 7648
rect 5021 7584 5027 7648
rect 4711 7583 5027 7584
rect 6781 7648 7097 7649
rect 6781 7584 6787 7648
rect 6851 7584 6867 7648
rect 6931 7584 6947 7648
rect 7011 7584 7027 7648
rect 7091 7584 7097 7648
rect 6781 7583 7097 7584
rect 8851 7648 9167 7649
rect 8851 7584 8857 7648
rect 8921 7584 8937 7648
rect 9001 7584 9017 7648
rect 9081 7584 9097 7648
rect 9161 7584 9167 7648
rect 8851 7583 9167 7584
rect 1981 7104 2297 7105
rect 1981 7040 1987 7104
rect 2051 7040 2067 7104
rect 2131 7040 2147 7104
rect 2211 7040 2227 7104
rect 2291 7040 2297 7104
rect 1981 7039 2297 7040
rect 4051 7104 4367 7105
rect 4051 7040 4057 7104
rect 4121 7040 4137 7104
rect 4201 7040 4217 7104
rect 4281 7040 4297 7104
rect 4361 7040 4367 7104
rect 4051 7039 4367 7040
rect 6121 7104 6437 7105
rect 6121 7040 6127 7104
rect 6191 7040 6207 7104
rect 6271 7040 6287 7104
rect 6351 7040 6367 7104
rect 6431 7040 6437 7104
rect 6121 7039 6437 7040
rect 8191 7104 8507 7105
rect 8191 7040 8197 7104
rect 8261 7040 8277 7104
rect 8341 7040 8357 7104
rect 8421 7040 8437 7104
rect 8501 7040 8507 7104
rect 8191 7039 8507 7040
rect 0 6898 800 6928
rect 1485 6898 1551 6901
rect 0 6896 1551 6898
rect 0 6840 1490 6896
rect 1546 6840 1551 6896
rect 0 6838 1551 6840
rect 0 6808 800 6838
rect 1485 6835 1551 6838
rect 2641 6560 2957 6561
rect 2641 6496 2647 6560
rect 2711 6496 2727 6560
rect 2791 6496 2807 6560
rect 2871 6496 2887 6560
rect 2951 6496 2957 6560
rect 2641 6495 2957 6496
rect 4711 6560 5027 6561
rect 4711 6496 4717 6560
rect 4781 6496 4797 6560
rect 4861 6496 4877 6560
rect 4941 6496 4957 6560
rect 5021 6496 5027 6560
rect 4711 6495 5027 6496
rect 6781 6560 7097 6561
rect 6781 6496 6787 6560
rect 6851 6496 6867 6560
rect 6931 6496 6947 6560
rect 7011 6496 7027 6560
rect 7091 6496 7097 6560
rect 6781 6495 7097 6496
rect 8851 6560 9167 6561
rect 8851 6496 8857 6560
rect 8921 6496 8937 6560
rect 9001 6496 9017 6560
rect 9081 6496 9097 6560
rect 9161 6496 9167 6560
rect 8851 6495 9167 6496
rect 8661 6218 8727 6221
rect 9767 6218 10567 6248
rect 8661 6216 10567 6218
rect 8661 6160 8666 6216
rect 8722 6160 10567 6216
rect 8661 6158 10567 6160
rect 8661 6155 8727 6158
rect 9767 6128 10567 6158
rect 1981 6016 2297 6017
rect 1981 5952 1987 6016
rect 2051 5952 2067 6016
rect 2131 5952 2147 6016
rect 2211 5952 2227 6016
rect 2291 5952 2297 6016
rect 1981 5951 2297 5952
rect 4051 6016 4367 6017
rect 4051 5952 4057 6016
rect 4121 5952 4137 6016
rect 4201 5952 4217 6016
rect 4281 5952 4297 6016
rect 4361 5952 4367 6016
rect 4051 5951 4367 5952
rect 6121 6016 6437 6017
rect 6121 5952 6127 6016
rect 6191 5952 6207 6016
rect 6271 5952 6287 6016
rect 6351 5952 6367 6016
rect 6431 5952 6437 6016
rect 6121 5951 6437 5952
rect 8191 6016 8507 6017
rect 8191 5952 8197 6016
rect 8261 5952 8277 6016
rect 8341 5952 8357 6016
rect 8421 5952 8437 6016
rect 8501 5952 8507 6016
rect 8191 5951 8507 5952
rect 2641 5472 2957 5473
rect 2641 5408 2647 5472
rect 2711 5408 2727 5472
rect 2791 5408 2807 5472
rect 2871 5408 2887 5472
rect 2951 5408 2957 5472
rect 2641 5407 2957 5408
rect 4711 5472 5027 5473
rect 4711 5408 4717 5472
rect 4781 5408 4797 5472
rect 4861 5408 4877 5472
rect 4941 5408 4957 5472
rect 5021 5408 5027 5472
rect 4711 5407 5027 5408
rect 6781 5472 7097 5473
rect 6781 5408 6787 5472
rect 6851 5408 6867 5472
rect 6931 5408 6947 5472
rect 7011 5408 7027 5472
rect 7091 5408 7097 5472
rect 6781 5407 7097 5408
rect 8851 5472 9167 5473
rect 8851 5408 8857 5472
rect 8921 5408 8937 5472
rect 9001 5408 9017 5472
rect 9081 5408 9097 5472
rect 9161 5408 9167 5472
rect 8851 5407 9167 5408
rect 1981 4928 2297 4929
rect 0 4858 800 4888
rect 1981 4864 1987 4928
rect 2051 4864 2067 4928
rect 2131 4864 2147 4928
rect 2211 4864 2227 4928
rect 2291 4864 2297 4928
rect 1981 4863 2297 4864
rect 4051 4928 4367 4929
rect 4051 4864 4057 4928
rect 4121 4864 4137 4928
rect 4201 4864 4217 4928
rect 4281 4864 4297 4928
rect 4361 4864 4367 4928
rect 4051 4863 4367 4864
rect 6121 4928 6437 4929
rect 6121 4864 6127 4928
rect 6191 4864 6207 4928
rect 6271 4864 6287 4928
rect 6351 4864 6367 4928
rect 6431 4864 6437 4928
rect 6121 4863 6437 4864
rect 8191 4928 8507 4929
rect 8191 4864 8197 4928
rect 8261 4864 8277 4928
rect 8341 4864 8357 4928
rect 8421 4864 8437 4928
rect 8501 4864 8507 4928
rect 8191 4863 8507 4864
rect 933 4858 999 4861
rect 0 4856 999 4858
rect 0 4800 938 4856
rect 994 4800 999 4856
rect 0 4798 999 4800
rect 0 4768 800 4798
rect 933 4795 999 4798
rect 9029 4858 9095 4861
rect 9767 4858 10567 4888
rect 9029 4856 10567 4858
rect 9029 4800 9034 4856
rect 9090 4800 10567 4856
rect 9029 4798 10567 4800
rect 9029 4795 9095 4798
rect 9767 4768 10567 4798
rect 2641 4384 2957 4385
rect 2641 4320 2647 4384
rect 2711 4320 2727 4384
rect 2791 4320 2807 4384
rect 2871 4320 2887 4384
rect 2951 4320 2957 4384
rect 2641 4319 2957 4320
rect 4711 4384 5027 4385
rect 4711 4320 4717 4384
rect 4781 4320 4797 4384
rect 4861 4320 4877 4384
rect 4941 4320 4957 4384
rect 5021 4320 5027 4384
rect 4711 4319 5027 4320
rect 6781 4384 7097 4385
rect 6781 4320 6787 4384
rect 6851 4320 6867 4384
rect 6931 4320 6947 4384
rect 7011 4320 7027 4384
rect 7091 4320 7097 4384
rect 6781 4319 7097 4320
rect 8851 4384 9167 4385
rect 8851 4320 8857 4384
rect 8921 4320 8937 4384
rect 9001 4320 9017 4384
rect 9081 4320 9097 4384
rect 9161 4320 9167 4384
rect 8851 4319 9167 4320
rect 1981 3840 2297 3841
rect 1981 3776 1987 3840
rect 2051 3776 2067 3840
rect 2131 3776 2147 3840
rect 2211 3776 2227 3840
rect 2291 3776 2297 3840
rect 1981 3775 2297 3776
rect 4051 3840 4367 3841
rect 4051 3776 4057 3840
rect 4121 3776 4137 3840
rect 4201 3776 4217 3840
rect 4281 3776 4297 3840
rect 4361 3776 4367 3840
rect 4051 3775 4367 3776
rect 6121 3840 6437 3841
rect 6121 3776 6127 3840
rect 6191 3776 6207 3840
rect 6271 3776 6287 3840
rect 6351 3776 6367 3840
rect 6431 3776 6437 3840
rect 6121 3775 6437 3776
rect 8191 3840 8507 3841
rect 8191 3776 8197 3840
rect 8261 3776 8277 3840
rect 8341 3776 8357 3840
rect 8421 3776 8437 3840
rect 8501 3776 8507 3840
rect 8191 3775 8507 3776
rect 0 3498 800 3528
rect 933 3498 999 3501
rect 0 3496 999 3498
rect 0 3440 938 3496
rect 994 3440 999 3496
rect 0 3438 999 3440
rect 0 3408 800 3438
rect 933 3435 999 3438
rect 2641 3296 2957 3297
rect 2641 3232 2647 3296
rect 2711 3232 2727 3296
rect 2791 3232 2807 3296
rect 2871 3232 2887 3296
rect 2951 3232 2957 3296
rect 2641 3231 2957 3232
rect 4711 3296 5027 3297
rect 4711 3232 4717 3296
rect 4781 3232 4797 3296
rect 4861 3232 4877 3296
rect 4941 3232 4957 3296
rect 5021 3232 5027 3296
rect 4711 3231 5027 3232
rect 6781 3296 7097 3297
rect 6781 3232 6787 3296
rect 6851 3232 6867 3296
rect 6931 3232 6947 3296
rect 7011 3232 7027 3296
rect 7091 3232 7097 3296
rect 6781 3231 7097 3232
rect 8851 3296 9167 3297
rect 8851 3232 8857 3296
rect 8921 3232 8937 3296
rect 9001 3232 9017 3296
rect 9081 3232 9097 3296
rect 9161 3232 9167 3296
rect 8851 3231 9167 3232
rect 9397 2818 9463 2821
rect 9767 2818 10567 2848
rect 9397 2816 10567 2818
rect 9397 2760 9402 2816
rect 9458 2760 10567 2816
rect 9397 2758 10567 2760
rect 9397 2755 9463 2758
rect 1981 2752 2297 2753
rect 1981 2688 1987 2752
rect 2051 2688 2067 2752
rect 2131 2688 2147 2752
rect 2211 2688 2227 2752
rect 2291 2688 2297 2752
rect 1981 2687 2297 2688
rect 4051 2752 4367 2753
rect 4051 2688 4057 2752
rect 4121 2688 4137 2752
rect 4201 2688 4217 2752
rect 4281 2688 4297 2752
rect 4361 2688 4367 2752
rect 4051 2687 4367 2688
rect 6121 2752 6437 2753
rect 6121 2688 6127 2752
rect 6191 2688 6207 2752
rect 6271 2688 6287 2752
rect 6351 2688 6367 2752
rect 6431 2688 6437 2752
rect 6121 2687 6437 2688
rect 8191 2752 8507 2753
rect 8191 2688 8197 2752
rect 8261 2688 8277 2752
rect 8341 2688 8357 2752
rect 8421 2688 8437 2752
rect 8501 2688 8507 2752
rect 9767 2728 10567 2758
rect 8191 2687 8507 2688
rect 2641 2208 2957 2209
rect 2641 2144 2647 2208
rect 2711 2144 2727 2208
rect 2791 2144 2807 2208
rect 2871 2144 2887 2208
rect 2951 2144 2957 2208
rect 2641 2143 2957 2144
rect 4711 2208 5027 2209
rect 4711 2144 4717 2208
rect 4781 2144 4797 2208
rect 4861 2144 4877 2208
rect 4941 2144 4957 2208
rect 5021 2144 5027 2208
rect 4711 2143 5027 2144
rect 6781 2208 7097 2209
rect 6781 2144 6787 2208
rect 6851 2144 6867 2208
rect 6931 2144 6947 2208
rect 7011 2144 7027 2208
rect 7091 2144 7097 2208
rect 6781 2143 7097 2144
rect 8851 2208 9167 2209
rect 8851 2144 8857 2208
rect 8921 2144 8937 2208
rect 9001 2144 9017 2208
rect 9081 2144 9097 2208
rect 9161 2144 9167 2208
rect 8851 2143 9167 2144
rect 0 1458 800 1488
rect 1209 1458 1275 1461
rect 0 1456 1275 1458
rect 0 1400 1214 1456
rect 1270 1400 1275 1456
rect 0 1398 1275 1400
rect 0 1368 800 1398
rect 1209 1395 1275 1398
rect 8017 778 8083 781
rect 9767 778 10567 808
rect 8017 776 10567 778
rect 8017 720 8022 776
rect 8078 720 10567 776
rect 8017 718 10567 720
rect 8017 715 8083 718
rect 9767 688 10567 718
<< via3 >>
rect 1987 10364 2051 10368
rect 1987 10308 1991 10364
rect 1991 10308 2047 10364
rect 2047 10308 2051 10364
rect 1987 10304 2051 10308
rect 2067 10364 2131 10368
rect 2067 10308 2071 10364
rect 2071 10308 2127 10364
rect 2127 10308 2131 10364
rect 2067 10304 2131 10308
rect 2147 10364 2211 10368
rect 2147 10308 2151 10364
rect 2151 10308 2207 10364
rect 2207 10308 2211 10364
rect 2147 10304 2211 10308
rect 2227 10364 2291 10368
rect 2227 10308 2231 10364
rect 2231 10308 2287 10364
rect 2287 10308 2291 10364
rect 2227 10304 2291 10308
rect 4057 10364 4121 10368
rect 4057 10308 4061 10364
rect 4061 10308 4117 10364
rect 4117 10308 4121 10364
rect 4057 10304 4121 10308
rect 4137 10364 4201 10368
rect 4137 10308 4141 10364
rect 4141 10308 4197 10364
rect 4197 10308 4201 10364
rect 4137 10304 4201 10308
rect 4217 10364 4281 10368
rect 4217 10308 4221 10364
rect 4221 10308 4277 10364
rect 4277 10308 4281 10364
rect 4217 10304 4281 10308
rect 4297 10364 4361 10368
rect 4297 10308 4301 10364
rect 4301 10308 4357 10364
rect 4357 10308 4361 10364
rect 4297 10304 4361 10308
rect 6127 10364 6191 10368
rect 6127 10308 6131 10364
rect 6131 10308 6187 10364
rect 6187 10308 6191 10364
rect 6127 10304 6191 10308
rect 6207 10364 6271 10368
rect 6207 10308 6211 10364
rect 6211 10308 6267 10364
rect 6267 10308 6271 10364
rect 6207 10304 6271 10308
rect 6287 10364 6351 10368
rect 6287 10308 6291 10364
rect 6291 10308 6347 10364
rect 6347 10308 6351 10364
rect 6287 10304 6351 10308
rect 6367 10364 6431 10368
rect 6367 10308 6371 10364
rect 6371 10308 6427 10364
rect 6427 10308 6431 10364
rect 6367 10304 6431 10308
rect 8197 10364 8261 10368
rect 8197 10308 8201 10364
rect 8201 10308 8257 10364
rect 8257 10308 8261 10364
rect 8197 10304 8261 10308
rect 8277 10364 8341 10368
rect 8277 10308 8281 10364
rect 8281 10308 8337 10364
rect 8337 10308 8341 10364
rect 8277 10304 8341 10308
rect 8357 10364 8421 10368
rect 8357 10308 8361 10364
rect 8361 10308 8417 10364
rect 8417 10308 8421 10364
rect 8357 10304 8421 10308
rect 8437 10364 8501 10368
rect 8437 10308 8441 10364
rect 8441 10308 8497 10364
rect 8497 10308 8501 10364
rect 8437 10304 8501 10308
rect 2647 9820 2711 9824
rect 2647 9764 2651 9820
rect 2651 9764 2707 9820
rect 2707 9764 2711 9820
rect 2647 9760 2711 9764
rect 2727 9820 2791 9824
rect 2727 9764 2731 9820
rect 2731 9764 2787 9820
rect 2787 9764 2791 9820
rect 2727 9760 2791 9764
rect 2807 9820 2871 9824
rect 2807 9764 2811 9820
rect 2811 9764 2867 9820
rect 2867 9764 2871 9820
rect 2807 9760 2871 9764
rect 2887 9820 2951 9824
rect 2887 9764 2891 9820
rect 2891 9764 2947 9820
rect 2947 9764 2951 9820
rect 2887 9760 2951 9764
rect 4717 9820 4781 9824
rect 4717 9764 4721 9820
rect 4721 9764 4777 9820
rect 4777 9764 4781 9820
rect 4717 9760 4781 9764
rect 4797 9820 4861 9824
rect 4797 9764 4801 9820
rect 4801 9764 4857 9820
rect 4857 9764 4861 9820
rect 4797 9760 4861 9764
rect 4877 9820 4941 9824
rect 4877 9764 4881 9820
rect 4881 9764 4937 9820
rect 4937 9764 4941 9820
rect 4877 9760 4941 9764
rect 4957 9820 5021 9824
rect 4957 9764 4961 9820
rect 4961 9764 5017 9820
rect 5017 9764 5021 9820
rect 4957 9760 5021 9764
rect 6787 9820 6851 9824
rect 6787 9764 6791 9820
rect 6791 9764 6847 9820
rect 6847 9764 6851 9820
rect 6787 9760 6851 9764
rect 6867 9820 6931 9824
rect 6867 9764 6871 9820
rect 6871 9764 6927 9820
rect 6927 9764 6931 9820
rect 6867 9760 6931 9764
rect 6947 9820 7011 9824
rect 6947 9764 6951 9820
rect 6951 9764 7007 9820
rect 7007 9764 7011 9820
rect 6947 9760 7011 9764
rect 7027 9820 7091 9824
rect 7027 9764 7031 9820
rect 7031 9764 7087 9820
rect 7087 9764 7091 9820
rect 7027 9760 7091 9764
rect 8857 9820 8921 9824
rect 8857 9764 8861 9820
rect 8861 9764 8917 9820
rect 8917 9764 8921 9820
rect 8857 9760 8921 9764
rect 8937 9820 9001 9824
rect 8937 9764 8941 9820
rect 8941 9764 8997 9820
rect 8997 9764 9001 9820
rect 8937 9760 9001 9764
rect 9017 9820 9081 9824
rect 9017 9764 9021 9820
rect 9021 9764 9077 9820
rect 9077 9764 9081 9820
rect 9017 9760 9081 9764
rect 9097 9820 9161 9824
rect 9097 9764 9101 9820
rect 9101 9764 9157 9820
rect 9157 9764 9161 9820
rect 9097 9760 9161 9764
rect 1987 9276 2051 9280
rect 1987 9220 1991 9276
rect 1991 9220 2047 9276
rect 2047 9220 2051 9276
rect 1987 9216 2051 9220
rect 2067 9276 2131 9280
rect 2067 9220 2071 9276
rect 2071 9220 2127 9276
rect 2127 9220 2131 9276
rect 2067 9216 2131 9220
rect 2147 9276 2211 9280
rect 2147 9220 2151 9276
rect 2151 9220 2207 9276
rect 2207 9220 2211 9276
rect 2147 9216 2211 9220
rect 2227 9276 2291 9280
rect 2227 9220 2231 9276
rect 2231 9220 2287 9276
rect 2287 9220 2291 9276
rect 2227 9216 2291 9220
rect 4057 9276 4121 9280
rect 4057 9220 4061 9276
rect 4061 9220 4117 9276
rect 4117 9220 4121 9276
rect 4057 9216 4121 9220
rect 4137 9276 4201 9280
rect 4137 9220 4141 9276
rect 4141 9220 4197 9276
rect 4197 9220 4201 9276
rect 4137 9216 4201 9220
rect 4217 9276 4281 9280
rect 4217 9220 4221 9276
rect 4221 9220 4277 9276
rect 4277 9220 4281 9276
rect 4217 9216 4281 9220
rect 4297 9276 4361 9280
rect 4297 9220 4301 9276
rect 4301 9220 4357 9276
rect 4357 9220 4361 9276
rect 4297 9216 4361 9220
rect 6127 9276 6191 9280
rect 6127 9220 6131 9276
rect 6131 9220 6187 9276
rect 6187 9220 6191 9276
rect 6127 9216 6191 9220
rect 6207 9276 6271 9280
rect 6207 9220 6211 9276
rect 6211 9220 6267 9276
rect 6267 9220 6271 9276
rect 6207 9216 6271 9220
rect 6287 9276 6351 9280
rect 6287 9220 6291 9276
rect 6291 9220 6347 9276
rect 6347 9220 6351 9276
rect 6287 9216 6351 9220
rect 6367 9276 6431 9280
rect 6367 9220 6371 9276
rect 6371 9220 6427 9276
rect 6427 9220 6431 9276
rect 6367 9216 6431 9220
rect 8197 9276 8261 9280
rect 8197 9220 8201 9276
rect 8201 9220 8257 9276
rect 8257 9220 8261 9276
rect 8197 9216 8261 9220
rect 8277 9276 8341 9280
rect 8277 9220 8281 9276
rect 8281 9220 8337 9276
rect 8337 9220 8341 9276
rect 8277 9216 8341 9220
rect 8357 9276 8421 9280
rect 8357 9220 8361 9276
rect 8361 9220 8417 9276
rect 8417 9220 8421 9276
rect 8357 9216 8421 9220
rect 8437 9276 8501 9280
rect 8437 9220 8441 9276
rect 8441 9220 8497 9276
rect 8497 9220 8501 9276
rect 8437 9216 8501 9220
rect 2647 8732 2711 8736
rect 2647 8676 2651 8732
rect 2651 8676 2707 8732
rect 2707 8676 2711 8732
rect 2647 8672 2711 8676
rect 2727 8732 2791 8736
rect 2727 8676 2731 8732
rect 2731 8676 2787 8732
rect 2787 8676 2791 8732
rect 2727 8672 2791 8676
rect 2807 8732 2871 8736
rect 2807 8676 2811 8732
rect 2811 8676 2867 8732
rect 2867 8676 2871 8732
rect 2807 8672 2871 8676
rect 2887 8732 2951 8736
rect 2887 8676 2891 8732
rect 2891 8676 2947 8732
rect 2947 8676 2951 8732
rect 2887 8672 2951 8676
rect 4717 8732 4781 8736
rect 4717 8676 4721 8732
rect 4721 8676 4777 8732
rect 4777 8676 4781 8732
rect 4717 8672 4781 8676
rect 4797 8732 4861 8736
rect 4797 8676 4801 8732
rect 4801 8676 4857 8732
rect 4857 8676 4861 8732
rect 4797 8672 4861 8676
rect 4877 8732 4941 8736
rect 4877 8676 4881 8732
rect 4881 8676 4937 8732
rect 4937 8676 4941 8732
rect 4877 8672 4941 8676
rect 4957 8732 5021 8736
rect 4957 8676 4961 8732
rect 4961 8676 5017 8732
rect 5017 8676 5021 8732
rect 4957 8672 5021 8676
rect 6787 8732 6851 8736
rect 6787 8676 6791 8732
rect 6791 8676 6847 8732
rect 6847 8676 6851 8732
rect 6787 8672 6851 8676
rect 6867 8732 6931 8736
rect 6867 8676 6871 8732
rect 6871 8676 6927 8732
rect 6927 8676 6931 8732
rect 6867 8672 6931 8676
rect 6947 8732 7011 8736
rect 6947 8676 6951 8732
rect 6951 8676 7007 8732
rect 7007 8676 7011 8732
rect 6947 8672 7011 8676
rect 7027 8732 7091 8736
rect 7027 8676 7031 8732
rect 7031 8676 7087 8732
rect 7087 8676 7091 8732
rect 7027 8672 7091 8676
rect 8857 8732 8921 8736
rect 8857 8676 8861 8732
rect 8861 8676 8917 8732
rect 8917 8676 8921 8732
rect 8857 8672 8921 8676
rect 8937 8732 9001 8736
rect 8937 8676 8941 8732
rect 8941 8676 8997 8732
rect 8997 8676 9001 8732
rect 8937 8672 9001 8676
rect 9017 8732 9081 8736
rect 9017 8676 9021 8732
rect 9021 8676 9077 8732
rect 9077 8676 9081 8732
rect 9017 8672 9081 8676
rect 9097 8732 9161 8736
rect 9097 8676 9101 8732
rect 9101 8676 9157 8732
rect 9157 8676 9161 8732
rect 9097 8672 9161 8676
rect 1987 8188 2051 8192
rect 1987 8132 1991 8188
rect 1991 8132 2047 8188
rect 2047 8132 2051 8188
rect 1987 8128 2051 8132
rect 2067 8188 2131 8192
rect 2067 8132 2071 8188
rect 2071 8132 2127 8188
rect 2127 8132 2131 8188
rect 2067 8128 2131 8132
rect 2147 8188 2211 8192
rect 2147 8132 2151 8188
rect 2151 8132 2207 8188
rect 2207 8132 2211 8188
rect 2147 8128 2211 8132
rect 2227 8188 2291 8192
rect 2227 8132 2231 8188
rect 2231 8132 2287 8188
rect 2287 8132 2291 8188
rect 2227 8128 2291 8132
rect 4057 8188 4121 8192
rect 4057 8132 4061 8188
rect 4061 8132 4117 8188
rect 4117 8132 4121 8188
rect 4057 8128 4121 8132
rect 4137 8188 4201 8192
rect 4137 8132 4141 8188
rect 4141 8132 4197 8188
rect 4197 8132 4201 8188
rect 4137 8128 4201 8132
rect 4217 8188 4281 8192
rect 4217 8132 4221 8188
rect 4221 8132 4277 8188
rect 4277 8132 4281 8188
rect 4217 8128 4281 8132
rect 4297 8188 4361 8192
rect 4297 8132 4301 8188
rect 4301 8132 4357 8188
rect 4357 8132 4361 8188
rect 4297 8128 4361 8132
rect 6127 8188 6191 8192
rect 6127 8132 6131 8188
rect 6131 8132 6187 8188
rect 6187 8132 6191 8188
rect 6127 8128 6191 8132
rect 6207 8188 6271 8192
rect 6207 8132 6211 8188
rect 6211 8132 6267 8188
rect 6267 8132 6271 8188
rect 6207 8128 6271 8132
rect 6287 8188 6351 8192
rect 6287 8132 6291 8188
rect 6291 8132 6347 8188
rect 6347 8132 6351 8188
rect 6287 8128 6351 8132
rect 6367 8188 6431 8192
rect 6367 8132 6371 8188
rect 6371 8132 6427 8188
rect 6427 8132 6431 8188
rect 6367 8128 6431 8132
rect 8197 8188 8261 8192
rect 8197 8132 8201 8188
rect 8201 8132 8257 8188
rect 8257 8132 8261 8188
rect 8197 8128 8261 8132
rect 8277 8188 8341 8192
rect 8277 8132 8281 8188
rect 8281 8132 8337 8188
rect 8337 8132 8341 8188
rect 8277 8128 8341 8132
rect 8357 8188 8421 8192
rect 8357 8132 8361 8188
rect 8361 8132 8417 8188
rect 8417 8132 8421 8188
rect 8357 8128 8421 8132
rect 8437 8188 8501 8192
rect 8437 8132 8441 8188
rect 8441 8132 8497 8188
rect 8497 8132 8501 8188
rect 8437 8128 8501 8132
rect 2647 7644 2711 7648
rect 2647 7588 2651 7644
rect 2651 7588 2707 7644
rect 2707 7588 2711 7644
rect 2647 7584 2711 7588
rect 2727 7644 2791 7648
rect 2727 7588 2731 7644
rect 2731 7588 2787 7644
rect 2787 7588 2791 7644
rect 2727 7584 2791 7588
rect 2807 7644 2871 7648
rect 2807 7588 2811 7644
rect 2811 7588 2867 7644
rect 2867 7588 2871 7644
rect 2807 7584 2871 7588
rect 2887 7644 2951 7648
rect 2887 7588 2891 7644
rect 2891 7588 2947 7644
rect 2947 7588 2951 7644
rect 2887 7584 2951 7588
rect 4717 7644 4781 7648
rect 4717 7588 4721 7644
rect 4721 7588 4777 7644
rect 4777 7588 4781 7644
rect 4717 7584 4781 7588
rect 4797 7644 4861 7648
rect 4797 7588 4801 7644
rect 4801 7588 4857 7644
rect 4857 7588 4861 7644
rect 4797 7584 4861 7588
rect 4877 7644 4941 7648
rect 4877 7588 4881 7644
rect 4881 7588 4937 7644
rect 4937 7588 4941 7644
rect 4877 7584 4941 7588
rect 4957 7644 5021 7648
rect 4957 7588 4961 7644
rect 4961 7588 5017 7644
rect 5017 7588 5021 7644
rect 4957 7584 5021 7588
rect 6787 7644 6851 7648
rect 6787 7588 6791 7644
rect 6791 7588 6847 7644
rect 6847 7588 6851 7644
rect 6787 7584 6851 7588
rect 6867 7644 6931 7648
rect 6867 7588 6871 7644
rect 6871 7588 6927 7644
rect 6927 7588 6931 7644
rect 6867 7584 6931 7588
rect 6947 7644 7011 7648
rect 6947 7588 6951 7644
rect 6951 7588 7007 7644
rect 7007 7588 7011 7644
rect 6947 7584 7011 7588
rect 7027 7644 7091 7648
rect 7027 7588 7031 7644
rect 7031 7588 7087 7644
rect 7087 7588 7091 7644
rect 7027 7584 7091 7588
rect 8857 7644 8921 7648
rect 8857 7588 8861 7644
rect 8861 7588 8917 7644
rect 8917 7588 8921 7644
rect 8857 7584 8921 7588
rect 8937 7644 9001 7648
rect 8937 7588 8941 7644
rect 8941 7588 8997 7644
rect 8997 7588 9001 7644
rect 8937 7584 9001 7588
rect 9017 7644 9081 7648
rect 9017 7588 9021 7644
rect 9021 7588 9077 7644
rect 9077 7588 9081 7644
rect 9017 7584 9081 7588
rect 9097 7644 9161 7648
rect 9097 7588 9101 7644
rect 9101 7588 9157 7644
rect 9157 7588 9161 7644
rect 9097 7584 9161 7588
rect 1987 7100 2051 7104
rect 1987 7044 1991 7100
rect 1991 7044 2047 7100
rect 2047 7044 2051 7100
rect 1987 7040 2051 7044
rect 2067 7100 2131 7104
rect 2067 7044 2071 7100
rect 2071 7044 2127 7100
rect 2127 7044 2131 7100
rect 2067 7040 2131 7044
rect 2147 7100 2211 7104
rect 2147 7044 2151 7100
rect 2151 7044 2207 7100
rect 2207 7044 2211 7100
rect 2147 7040 2211 7044
rect 2227 7100 2291 7104
rect 2227 7044 2231 7100
rect 2231 7044 2287 7100
rect 2287 7044 2291 7100
rect 2227 7040 2291 7044
rect 4057 7100 4121 7104
rect 4057 7044 4061 7100
rect 4061 7044 4117 7100
rect 4117 7044 4121 7100
rect 4057 7040 4121 7044
rect 4137 7100 4201 7104
rect 4137 7044 4141 7100
rect 4141 7044 4197 7100
rect 4197 7044 4201 7100
rect 4137 7040 4201 7044
rect 4217 7100 4281 7104
rect 4217 7044 4221 7100
rect 4221 7044 4277 7100
rect 4277 7044 4281 7100
rect 4217 7040 4281 7044
rect 4297 7100 4361 7104
rect 4297 7044 4301 7100
rect 4301 7044 4357 7100
rect 4357 7044 4361 7100
rect 4297 7040 4361 7044
rect 6127 7100 6191 7104
rect 6127 7044 6131 7100
rect 6131 7044 6187 7100
rect 6187 7044 6191 7100
rect 6127 7040 6191 7044
rect 6207 7100 6271 7104
rect 6207 7044 6211 7100
rect 6211 7044 6267 7100
rect 6267 7044 6271 7100
rect 6207 7040 6271 7044
rect 6287 7100 6351 7104
rect 6287 7044 6291 7100
rect 6291 7044 6347 7100
rect 6347 7044 6351 7100
rect 6287 7040 6351 7044
rect 6367 7100 6431 7104
rect 6367 7044 6371 7100
rect 6371 7044 6427 7100
rect 6427 7044 6431 7100
rect 6367 7040 6431 7044
rect 8197 7100 8261 7104
rect 8197 7044 8201 7100
rect 8201 7044 8257 7100
rect 8257 7044 8261 7100
rect 8197 7040 8261 7044
rect 8277 7100 8341 7104
rect 8277 7044 8281 7100
rect 8281 7044 8337 7100
rect 8337 7044 8341 7100
rect 8277 7040 8341 7044
rect 8357 7100 8421 7104
rect 8357 7044 8361 7100
rect 8361 7044 8417 7100
rect 8417 7044 8421 7100
rect 8357 7040 8421 7044
rect 8437 7100 8501 7104
rect 8437 7044 8441 7100
rect 8441 7044 8497 7100
rect 8497 7044 8501 7100
rect 8437 7040 8501 7044
rect 2647 6556 2711 6560
rect 2647 6500 2651 6556
rect 2651 6500 2707 6556
rect 2707 6500 2711 6556
rect 2647 6496 2711 6500
rect 2727 6556 2791 6560
rect 2727 6500 2731 6556
rect 2731 6500 2787 6556
rect 2787 6500 2791 6556
rect 2727 6496 2791 6500
rect 2807 6556 2871 6560
rect 2807 6500 2811 6556
rect 2811 6500 2867 6556
rect 2867 6500 2871 6556
rect 2807 6496 2871 6500
rect 2887 6556 2951 6560
rect 2887 6500 2891 6556
rect 2891 6500 2947 6556
rect 2947 6500 2951 6556
rect 2887 6496 2951 6500
rect 4717 6556 4781 6560
rect 4717 6500 4721 6556
rect 4721 6500 4777 6556
rect 4777 6500 4781 6556
rect 4717 6496 4781 6500
rect 4797 6556 4861 6560
rect 4797 6500 4801 6556
rect 4801 6500 4857 6556
rect 4857 6500 4861 6556
rect 4797 6496 4861 6500
rect 4877 6556 4941 6560
rect 4877 6500 4881 6556
rect 4881 6500 4937 6556
rect 4937 6500 4941 6556
rect 4877 6496 4941 6500
rect 4957 6556 5021 6560
rect 4957 6500 4961 6556
rect 4961 6500 5017 6556
rect 5017 6500 5021 6556
rect 4957 6496 5021 6500
rect 6787 6556 6851 6560
rect 6787 6500 6791 6556
rect 6791 6500 6847 6556
rect 6847 6500 6851 6556
rect 6787 6496 6851 6500
rect 6867 6556 6931 6560
rect 6867 6500 6871 6556
rect 6871 6500 6927 6556
rect 6927 6500 6931 6556
rect 6867 6496 6931 6500
rect 6947 6556 7011 6560
rect 6947 6500 6951 6556
rect 6951 6500 7007 6556
rect 7007 6500 7011 6556
rect 6947 6496 7011 6500
rect 7027 6556 7091 6560
rect 7027 6500 7031 6556
rect 7031 6500 7087 6556
rect 7087 6500 7091 6556
rect 7027 6496 7091 6500
rect 8857 6556 8921 6560
rect 8857 6500 8861 6556
rect 8861 6500 8917 6556
rect 8917 6500 8921 6556
rect 8857 6496 8921 6500
rect 8937 6556 9001 6560
rect 8937 6500 8941 6556
rect 8941 6500 8997 6556
rect 8997 6500 9001 6556
rect 8937 6496 9001 6500
rect 9017 6556 9081 6560
rect 9017 6500 9021 6556
rect 9021 6500 9077 6556
rect 9077 6500 9081 6556
rect 9017 6496 9081 6500
rect 9097 6556 9161 6560
rect 9097 6500 9101 6556
rect 9101 6500 9157 6556
rect 9157 6500 9161 6556
rect 9097 6496 9161 6500
rect 1987 6012 2051 6016
rect 1987 5956 1991 6012
rect 1991 5956 2047 6012
rect 2047 5956 2051 6012
rect 1987 5952 2051 5956
rect 2067 6012 2131 6016
rect 2067 5956 2071 6012
rect 2071 5956 2127 6012
rect 2127 5956 2131 6012
rect 2067 5952 2131 5956
rect 2147 6012 2211 6016
rect 2147 5956 2151 6012
rect 2151 5956 2207 6012
rect 2207 5956 2211 6012
rect 2147 5952 2211 5956
rect 2227 6012 2291 6016
rect 2227 5956 2231 6012
rect 2231 5956 2287 6012
rect 2287 5956 2291 6012
rect 2227 5952 2291 5956
rect 4057 6012 4121 6016
rect 4057 5956 4061 6012
rect 4061 5956 4117 6012
rect 4117 5956 4121 6012
rect 4057 5952 4121 5956
rect 4137 6012 4201 6016
rect 4137 5956 4141 6012
rect 4141 5956 4197 6012
rect 4197 5956 4201 6012
rect 4137 5952 4201 5956
rect 4217 6012 4281 6016
rect 4217 5956 4221 6012
rect 4221 5956 4277 6012
rect 4277 5956 4281 6012
rect 4217 5952 4281 5956
rect 4297 6012 4361 6016
rect 4297 5956 4301 6012
rect 4301 5956 4357 6012
rect 4357 5956 4361 6012
rect 4297 5952 4361 5956
rect 6127 6012 6191 6016
rect 6127 5956 6131 6012
rect 6131 5956 6187 6012
rect 6187 5956 6191 6012
rect 6127 5952 6191 5956
rect 6207 6012 6271 6016
rect 6207 5956 6211 6012
rect 6211 5956 6267 6012
rect 6267 5956 6271 6012
rect 6207 5952 6271 5956
rect 6287 6012 6351 6016
rect 6287 5956 6291 6012
rect 6291 5956 6347 6012
rect 6347 5956 6351 6012
rect 6287 5952 6351 5956
rect 6367 6012 6431 6016
rect 6367 5956 6371 6012
rect 6371 5956 6427 6012
rect 6427 5956 6431 6012
rect 6367 5952 6431 5956
rect 8197 6012 8261 6016
rect 8197 5956 8201 6012
rect 8201 5956 8257 6012
rect 8257 5956 8261 6012
rect 8197 5952 8261 5956
rect 8277 6012 8341 6016
rect 8277 5956 8281 6012
rect 8281 5956 8337 6012
rect 8337 5956 8341 6012
rect 8277 5952 8341 5956
rect 8357 6012 8421 6016
rect 8357 5956 8361 6012
rect 8361 5956 8417 6012
rect 8417 5956 8421 6012
rect 8357 5952 8421 5956
rect 8437 6012 8501 6016
rect 8437 5956 8441 6012
rect 8441 5956 8497 6012
rect 8497 5956 8501 6012
rect 8437 5952 8501 5956
rect 2647 5468 2711 5472
rect 2647 5412 2651 5468
rect 2651 5412 2707 5468
rect 2707 5412 2711 5468
rect 2647 5408 2711 5412
rect 2727 5468 2791 5472
rect 2727 5412 2731 5468
rect 2731 5412 2787 5468
rect 2787 5412 2791 5468
rect 2727 5408 2791 5412
rect 2807 5468 2871 5472
rect 2807 5412 2811 5468
rect 2811 5412 2867 5468
rect 2867 5412 2871 5468
rect 2807 5408 2871 5412
rect 2887 5468 2951 5472
rect 2887 5412 2891 5468
rect 2891 5412 2947 5468
rect 2947 5412 2951 5468
rect 2887 5408 2951 5412
rect 4717 5468 4781 5472
rect 4717 5412 4721 5468
rect 4721 5412 4777 5468
rect 4777 5412 4781 5468
rect 4717 5408 4781 5412
rect 4797 5468 4861 5472
rect 4797 5412 4801 5468
rect 4801 5412 4857 5468
rect 4857 5412 4861 5468
rect 4797 5408 4861 5412
rect 4877 5468 4941 5472
rect 4877 5412 4881 5468
rect 4881 5412 4937 5468
rect 4937 5412 4941 5468
rect 4877 5408 4941 5412
rect 4957 5468 5021 5472
rect 4957 5412 4961 5468
rect 4961 5412 5017 5468
rect 5017 5412 5021 5468
rect 4957 5408 5021 5412
rect 6787 5468 6851 5472
rect 6787 5412 6791 5468
rect 6791 5412 6847 5468
rect 6847 5412 6851 5468
rect 6787 5408 6851 5412
rect 6867 5468 6931 5472
rect 6867 5412 6871 5468
rect 6871 5412 6927 5468
rect 6927 5412 6931 5468
rect 6867 5408 6931 5412
rect 6947 5468 7011 5472
rect 6947 5412 6951 5468
rect 6951 5412 7007 5468
rect 7007 5412 7011 5468
rect 6947 5408 7011 5412
rect 7027 5468 7091 5472
rect 7027 5412 7031 5468
rect 7031 5412 7087 5468
rect 7087 5412 7091 5468
rect 7027 5408 7091 5412
rect 8857 5468 8921 5472
rect 8857 5412 8861 5468
rect 8861 5412 8917 5468
rect 8917 5412 8921 5468
rect 8857 5408 8921 5412
rect 8937 5468 9001 5472
rect 8937 5412 8941 5468
rect 8941 5412 8997 5468
rect 8997 5412 9001 5468
rect 8937 5408 9001 5412
rect 9017 5468 9081 5472
rect 9017 5412 9021 5468
rect 9021 5412 9077 5468
rect 9077 5412 9081 5468
rect 9017 5408 9081 5412
rect 9097 5468 9161 5472
rect 9097 5412 9101 5468
rect 9101 5412 9157 5468
rect 9157 5412 9161 5468
rect 9097 5408 9161 5412
rect 1987 4924 2051 4928
rect 1987 4868 1991 4924
rect 1991 4868 2047 4924
rect 2047 4868 2051 4924
rect 1987 4864 2051 4868
rect 2067 4924 2131 4928
rect 2067 4868 2071 4924
rect 2071 4868 2127 4924
rect 2127 4868 2131 4924
rect 2067 4864 2131 4868
rect 2147 4924 2211 4928
rect 2147 4868 2151 4924
rect 2151 4868 2207 4924
rect 2207 4868 2211 4924
rect 2147 4864 2211 4868
rect 2227 4924 2291 4928
rect 2227 4868 2231 4924
rect 2231 4868 2287 4924
rect 2287 4868 2291 4924
rect 2227 4864 2291 4868
rect 4057 4924 4121 4928
rect 4057 4868 4061 4924
rect 4061 4868 4117 4924
rect 4117 4868 4121 4924
rect 4057 4864 4121 4868
rect 4137 4924 4201 4928
rect 4137 4868 4141 4924
rect 4141 4868 4197 4924
rect 4197 4868 4201 4924
rect 4137 4864 4201 4868
rect 4217 4924 4281 4928
rect 4217 4868 4221 4924
rect 4221 4868 4277 4924
rect 4277 4868 4281 4924
rect 4217 4864 4281 4868
rect 4297 4924 4361 4928
rect 4297 4868 4301 4924
rect 4301 4868 4357 4924
rect 4357 4868 4361 4924
rect 4297 4864 4361 4868
rect 6127 4924 6191 4928
rect 6127 4868 6131 4924
rect 6131 4868 6187 4924
rect 6187 4868 6191 4924
rect 6127 4864 6191 4868
rect 6207 4924 6271 4928
rect 6207 4868 6211 4924
rect 6211 4868 6267 4924
rect 6267 4868 6271 4924
rect 6207 4864 6271 4868
rect 6287 4924 6351 4928
rect 6287 4868 6291 4924
rect 6291 4868 6347 4924
rect 6347 4868 6351 4924
rect 6287 4864 6351 4868
rect 6367 4924 6431 4928
rect 6367 4868 6371 4924
rect 6371 4868 6427 4924
rect 6427 4868 6431 4924
rect 6367 4864 6431 4868
rect 8197 4924 8261 4928
rect 8197 4868 8201 4924
rect 8201 4868 8257 4924
rect 8257 4868 8261 4924
rect 8197 4864 8261 4868
rect 8277 4924 8341 4928
rect 8277 4868 8281 4924
rect 8281 4868 8337 4924
rect 8337 4868 8341 4924
rect 8277 4864 8341 4868
rect 8357 4924 8421 4928
rect 8357 4868 8361 4924
rect 8361 4868 8417 4924
rect 8417 4868 8421 4924
rect 8357 4864 8421 4868
rect 8437 4924 8501 4928
rect 8437 4868 8441 4924
rect 8441 4868 8497 4924
rect 8497 4868 8501 4924
rect 8437 4864 8501 4868
rect 2647 4380 2711 4384
rect 2647 4324 2651 4380
rect 2651 4324 2707 4380
rect 2707 4324 2711 4380
rect 2647 4320 2711 4324
rect 2727 4380 2791 4384
rect 2727 4324 2731 4380
rect 2731 4324 2787 4380
rect 2787 4324 2791 4380
rect 2727 4320 2791 4324
rect 2807 4380 2871 4384
rect 2807 4324 2811 4380
rect 2811 4324 2867 4380
rect 2867 4324 2871 4380
rect 2807 4320 2871 4324
rect 2887 4380 2951 4384
rect 2887 4324 2891 4380
rect 2891 4324 2947 4380
rect 2947 4324 2951 4380
rect 2887 4320 2951 4324
rect 4717 4380 4781 4384
rect 4717 4324 4721 4380
rect 4721 4324 4777 4380
rect 4777 4324 4781 4380
rect 4717 4320 4781 4324
rect 4797 4380 4861 4384
rect 4797 4324 4801 4380
rect 4801 4324 4857 4380
rect 4857 4324 4861 4380
rect 4797 4320 4861 4324
rect 4877 4380 4941 4384
rect 4877 4324 4881 4380
rect 4881 4324 4937 4380
rect 4937 4324 4941 4380
rect 4877 4320 4941 4324
rect 4957 4380 5021 4384
rect 4957 4324 4961 4380
rect 4961 4324 5017 4380
rect 5017 4324 5021 4380
rect 4957 4320 5021 4324
rect 6787 4380 6851 4384
rect 6787 4324 6791 4380
rect 6791 4324 6847 4380
rect 6847 4324 6851 4380
rect 6787 4320 6851 4324
rect 6867 4380 6931 4384
rect 6867 4324 6871 4380
rect 6871 4324 6927 4380
rect 6927 4324 6931 4380
rect 6867 4320 6931 4324
rect 6947 4380 7011 4384
rect 6947 4324 6951 4380
rect 6951 4324 7007 4380
rect 7007 4324 7011 4380
rect 6947 4320 7011 4324
rect 7027 4380 7091 4384
rect 7027 4324 7031 4380
rect 7031 4324 7087 4380
rect 7087 4324 7091 4380
rect 7027 4320 7091 4324
rect 8857 4380 8921 4384
rect 8857 4324 8861 4380
rect 8861 4324 8917 4380
rect 8917 4324 8921 4380
rect 8857 4320 8921 4324
rect 8937 4380 9001 4384
rect 8937 4324 8941 4380
rect 8941 4324 8997 4380
rect 8997 4324 9001 4380
rect 8937 4320 9001 4324
rect 9017 4380 9081 4384
rect 9017 4324 9021 4380
rect 9021 4324 9077 4380
rect 9077 4324 9081 4380
rect 9017 4320 9081 4324
rect 9097 4380 9161 4384
rect 9097 4324 9101 4380
rect 9101 4324 9157 4380
rect 9157 4324 9161 4380
rect 9097 4320 9161 4324
rect 1987 3836 2051 3840
rect 1987 3780 1991 3836
rect 1991 3780 2047 3836
rect 2047 3780 2051 3836
rect 1987 3776 2051 3780
rect 2067 3836 2131 3840
rect 2067 3780 2071 3836
rect 2071 3780 2127 3836
rect 2127 3780 2131 3836
rect 2067 3776 2131 3780
rect 2147 3836 2211 3840
rect 2147 3780 2151 3836
rect 2151 3780 2207 3836
rect 2207 3780 2211 3836
rect 2147 3776 2211 3780
rect 2227 3836 2291 3840
rect 2227 3780 2231 3836
rect 2231 3780 2287 3836
rect 2287 3780 2291 3836
rect 2227 3776 2291 3780
rect 4057 3836 4121 3840
rect 4057 3780 4061 3836
rect 4061 3780 4117 3836
rect 4117 3780 4121 3836
rect 4057 3776 4121 3780
rect 4137 3836 4201 3840
rect 4137 3780 4141 3836
rect 4141 3780 4197 3836
rect 4197 3780 4201 3836
rect 4137 3776 4201 3780
rect 4217 3836 4281 3840
rect 4217 3780 4221 3836
rect 4221 3780 4277 3836
rect 4277 3780 4281 3836
rect 4217 3776 4281 3780
rect 4297 3836 4361 3840
rect 4297 3780 4301 3836
rect 4301 3780 4357 3836
rect 4357 3780 4361 3836
rect 4297 3776 4361 3780
rect 6127 3836 6191 3840
rect 6127 3780 6131 3836
rect 6131 3780 6187 3836
rect 6187 3780 6191 3836
rect 6127 3776 6191 3780
rect 6207 3836 6271 3840
rect 6207 3780 6211 3836
rect 6211 3780 6267 3836
rect 6267 3780 6271 3836
rect 6207 3776 6271 3780
rect 6287 3836 6351 3840
rect 6287 3780 6291 3836
rect 6291 3780 6347 3836
rect 6347 3780 6351 3836
rect 6287 3776 6351 3780
rect 6367 3836 6431 3840
rect 6367 3780 6371 3836
rect 6371 3780 6427 3836
rect 6427 3780 6431 3836
rect 6367 3776 6431 3780
rect 8197 3836 8261 3840
rect 8197 3780 8201 3836
rect 8201 3780 8257 3836
rect 8257 3780 8261 3836
rect 8197 3776 8261 3780
rect 8277 3836 8341 3840
rect 8277 3780 8281 3836
rect 8281 3780 8337 3836
rect 8337 3780 8341 3836
rect 8277 3776 8341 3780
rect 8357 3836 8421 3840
rect 8357 3780 8361 3836
rect 8361 3780 8417 3836
rect 8417 3780 8421 3836
rect 8357 3776 8421 3780
rect 8437 3836 8501 3840
rect 8437 3780 8441 3836
rect 8441 3780 8497 3836
rect 8497 3780 8501 3836
rect 8437 3776 8501 3780
rect 2647 3292 2711 3296
rect 2647 3236 2651 3292
rect 2651 3236 2707 3292
rect 2707 3236 2711 3292
rect 2647 3232 2711 3236
rect 2727 3292 2791 3296
rect 2727 3236 2731 3292
rect 2731 3236 2787 3292
rect 2787 3236 2791 3292
rect 2727 3232 2791 3236
rect 2807 3292 2871 3296
rect 2807 3236 2811 3292
rect 2811 3236 2867 3292
rect 2867 3236 2871 3292
rect 2807 3232 2871 3236
rect 2887 3292 2951 3296
rect 2887 3236 2891 3292
rect 2891 3236 2947 3292
rect 2947 3236 2951 3292
rect 2887 3232 2951 3236
rect 4717 3292 4781 3296
rect 4717 3236 4721 3292
rect 4721 3236 4777 3292
rect 4777 3236 4781 3292
rect 4717 3232 4781 3236
rect 4797 3292 4861 3296
rect 4797 3236 4801 3292
rect 4801 3236 4857 3292
rect 4857 3236 4861 3292
rect 4797 3232 4861 3236
rect 4877 3292 4941 3296
rect 4877 3236 4881 3292
rect 4881 3236 4937 3292
rect 4937 3236 4941 3292
rect 4877 3232 4941 3236
rect 4957 3292 5021 3296
rect 4957 3236 4961 3292
rect 4961 3236 5017 3292
rect 5017 3236 5021 3292
rect 4957 3232 5021 3236
rect 6787 3292 6851 3296
rect 6787 3236 6791 3292
rect 6791 3236 6847 3292
rect 6847 3236 6851 3292
rect 6787 3232 6851 3236
rect 6867 3292 6931 3296
rect 6867 3236 6871 3292
rect 6871 3236 6927 3292
rect 6927 3236 6931 3292
rect 6867 3232 6931 3236
rect 6947 3292 7011 3296
rect 6947 3236 6951 3292
rect 6951 3236 7007 3292
rect 7007 3236 7011 3292
rect 6947 3232 7011 3236
rect 7027 3292 7091 3296
rect 7027 3236 7031 3292
rect 7031 3236 7087 3292
rect 7087 3236 7091 3292
rect 7027 3232 7091 3236
rect 8857 3292 8921 3296
rect 8857 3236 8861 3292
rect 8861 3236 8917 3292
rect 8917 3236 8921 3292
rect 8857 3232 8921 3236
rect 8937 3292 9001 3296
rect 8937 3236 8941 3292
rect 8941 3236 8997 3292
rect 8997 3236 9001 3292
rect 8937 3232 9001 3236
rect 9017 3292 9081 3296
rect 9017 3236 9021 3292
rect 9021 3236 9077 3292
rect 9077 3236 9081 3292
rect 9017 3232 9081 3236
rect 9097 3292 9161 3296
rect 9097 3236 9101 3292
rect 9101 3236 9157 3292
rect 9157 3236 9161 3292
rect 9097 3232 9161 3236
rect 1987 2748 2051 2752
rect 1987 2692 1991 2748
rect 1991 2692 2047 2748
rect 2047 2692 2051 2748
rect 1987 2688 2051 2692
rect 2067 2748 2131 2752
rect 2067 2692 2071 2748
rect 2071 2692 2127 2748
rect 2127 2692 2131 2748
rect 2067 2688 2131 2692
rect 2147 2748 2211 2752
rect 2147 2692 2151 2748
rect 2151 2692 2207 2748
rect 2207 2692 2211 2748
rect 2147 2688 2211 2692
rect 2227 2748 2291 2752
rect 2227 2692 2231 2748
rect 2231 2692 2287 2748
rect 2287 2692 2291 2748
rect 2227 2688 2291 2692
rect 4057 2748 4121 2752
rect 4057 2692 4061 2748
rect 4061 2692 4117 2748
rect 4117 2692 4121 2748
rect 4057 2688 4121 2692
rect 4137 2748 4201 2752
rect 4137 2692 4141 2748
rect 4141 2692 4197 2748
rect 4197 2692 4201 2748
rect 4137 2688 4201 2692
rect 4217 2748 4281 2752
rect 4217 2692 4221 2748
rect 4221 2692 4277 2748
rect 4277 2692 4281 2748
rect 4217 2688 4281 2692
rect 4297 2748 4361 2752
rect 4297 2692 4301 2748
rect 4301 2692 4357 2748
rect 4357 2692 4361 2748
rect 4297 2688 4361 2692
rect 6127 2748 6191 2752
rect 6127 2692 6131 2748
rect 6131 2692 6187 2748
rect 6187 2692 6191 2748
rect 6127 2688 6191 2692
rect 6207 2748 6271 2752
rect 6207 2692 6211 2748
rect 6211 2692 6267 2748
rect 6267 2692 6271 2748
rect 6207 2688 6271 2692
rect 6287 2748 6351 2752
rect 6287 2692 6291 2748
rect 6291 2692 6347 2748
rect 6347 2692 6351 2748
rect 6287 2688 6351 2692
rect 6367 2748 6431 2752
rect 6367 2692 6371 2748
rect 6371 2692 6427 2748
rect 6427 2692 6431 2748
rect 6367 2688 6431 2692
rect 8197 2748 8261 2752
rect 8197 2692 8201 2748
rect 8201 2692 8257 2748
rect 8257 2692 8261 2748
rect 8197 2688 8261 2692
rect 8277 2748 8341 2752
rect 8277 2692 8281 2748
rect 8281 2692 8337 2748
rect 8337 2692 8341 2748
rect 8277 2688 8341 2692
rect 8357 2748 8421 2752
rect 8357 2692 8361 2748
rect 8361 2692 8417 2748
rect 8417 2692 8421 2748
rect 8357 2688 8421 2692
rect 8437 2748 8501 2752
rect 8437 2692 8441 2748
rect 8441 2692 8497 2748
rect 8497 2692 8501 2748
rect 8437 2688 8501 2692
rect 2647 2204 2711 2208
rect 2647 2148 2651 2204
rect 2651 2148 2707 2204
rect 2707 2148 2711 2204
rect 2647 2144 2711 2148
rect 2727 2204 2791 2208
rect 2727 2148 2731 2204
rect 2731 2148 2787 2204
rect 2787 2148 2791 2204
rect 2727 2144 2791 2148
rect 2807 2204 2871 2208
rect 2807 2148 2811 2204
rect 2811 2148 2867 2204
rect 2867 2148 2871 2204
rect 2807 2144 2871 2148
rect 2887 2204 2951 2208
rect 2887 2148 2891 2204
rect 2891 2148 2947 2204
rect 2947 2148 2951 2204
rect 2887 2144 2951 2148
rect 4717 2204 4781 2208
rect 4717 2148 4721 2204
rect 4721 2148 4777 2204
rect 4777 2148 4781 2204
rect 4717 2144 4781 2148
rect 4797 2204 4861 2208
rect 4797 2148 4801 2204
rect 4801 2148 4857 2204
rect 4857 2148 4861 2204
rect 4797 2144 4861 2148
rect 4877 2204 4941 2208
rect 4877 2148 4881 2204
rect 4881 2148 4937 2204
rect 4937 2148 4941 2204
rect 4877 2144 4941 2148
rect 4957 2204 5021 2208
rect 4957 2148 4961 2204
rect 4961 2148 5017 2204
rect 5017 2148 5021 2204
rect 4957 2144 5021 2148
rect 6787 2204 6851 2208
rect 6787 2148 6791 2204
rect 6791 2148 6847 2204
rect 6847 2148 6851 2204
rect 6787 2144 6851 2148
rect 6867 2204 6931 2208
rect 6867 2148 6871 2204
rect 6871 2148 6927 2204
rect 6927 2148 6931 2204
rect 6867 2144 6931 2148
rect 6947 2204 7011 2208
rect 6947 2148 6951 2204
rect 6951 2148 7007 2204
rect 7007 2148 7011 2204
rect 6947 2144 7011 2148
rect 7027 2204 7091 2208
rect 7027 2148 7031 2204
rect 7031 2148 7087 2204
rect 7087 2148 7091 2204
rect 7027 2144 7091 2148
rect 8857 2204 8921 2208
rect 8857 2148 8861 2204
rect 8861 2148 8917 2204
rect 8917 2148 8921 2204
rect 8857 2144 8921 2148
rect 8937 2204 9001 2208
rect 8937 2148 8941 2204
rect 8941 2148 8997 2204
rect 8997 2148 9001 2204
rect 8937 2144 9001 2148
rect 9017 2204 9081 2208
rect 9017 2148 9021 2204
rect 9021 2148 9077 2204
rect 9077 2148 9081 2204
rect 9017 2144 9081 2148
rect 9097 2204 9161 2208
rect 9097 2148 9101 2204
rect 9101 2148 9157 2204
rect 9157 2148 9161 2204
rect 9097 2144 9161 2148
<< metal4 >>
rect 1979 10368 2299 10384
rect 1979 10304 1987 10368
rect 2051 10304 2067 10368
rect 2131 10304 2147 10368
rect 2211 10304 2227 10368
rect 2291 10304 2299 10368
rect 1979 9434 2299 10304
rect 1979 9280 2021 9434
rect 2257 9280 2299 9434
rect 1979 9216 1987 9280
rect 2291 9216 2299 9280
rect 1979 9198 2021 9216
rect 2257 9198 2299 9216
rect 1979 8192 2299 9198
rect 1979 8128 1987 8192
rect 2051 8128 2067 8192
rect 2131 8128 2147 8192
rect 2211 8128 2227 8192
rect 2291 8128 2299 8192
rect 1979 7394 2299 8128
rect 1979 7158 2021 7394
rect 2257 7158 2299 7394
rect 1979 7104 2299 7158
rect 1979 7040 1987 7104
rect 2051 7040 2067 7104
rect 2131 7040 2147 7104
rect 2211 7040 2227 7104
rect 2291 7040 2299 7104
rect 1979 6016 2299 7040
rect 1979 5952 1987 6016
rect 2051 5952 2067 6016
rect 2131 5952 2147 6016
rect 2211 5952 2227 6016
rect 2291 5952 2299 6016
rect 1979 5354 2299 5952
rect 1979 5118 2021 5354
rect 2257 5118 2299 5354
rect 1979 4928 2299 5118
rect 1979 4864 1987 4928
rect 2051 4864 2067 4928
rect 2131 4864 2147 4928
rect 2211 4864 2227 4928
rect 2291 4864 2299 4928
rect 1979 3840 2299 4864
rect 1979 3776 1987 3840
rect 2051 3776 2067 3840
rect 2131 3776 2147 3840
rect 2211 3776 2227 3840
rect 2291 3776 2299 3840
rect 1979 3314 2299 3776
rect 1979 3078 2021 3314
rect 2257 3078 2299 3314
rect 1979 2752 2299 3078
rect 1979 2688 1987 2752
rect 2051 2688 2067 2752
rect 2131 2688 2147 2752
rect 2211 2688 2227 2752
rect 2291 2688 2299 2752
rect 1979 2128 2299 2688
rect 2639 10094 2959 10384
rect 2639 9858 2681 10094
rect 2917 9858 2959 10094
rect 2639 9824 2959 9858
rect 2639 9760 2647 9824
rect 2711 9760 2727 9824
rect 2791 9760 2807 9824
rect 2871 9760 2887 9824
rect 2951 9760 2959 9824
rect 2639 8736 2959 9760
rect 2639 8672 2647 8736
rect 2711 8672 2727 8736
rect 2791 8672 2807 8736
rect 2871 8672 2887 8736
rect 2951 8672 2959 8736
rect 2639 8054 2959 8672
rect 2639 7818 2681 8054
rect 2917 7818 2959 8054
rect 2639 7648 2959 7818
rect 2639 7584 2647 7648
rect 2711 7584 2727 7648
rect 2791 7584 2807 7648
rect 2871 7584 2887 7648
rect 2951 7584 2959 7648
rect 2639 6560 2959 7584
rect 2639 6496 2647 6560
rect 2711 6496 2727 6560
rect 2791 6496 2807 6560
rect 2871 6496 2887 6560
rect 2951 6496 2959 6560
rect 2639 6014 2959 6496
rect 2639 5778 2681 6014
rect 2917 5778 2959 6014
rect 2639 5472 2959 5778
rect 2639 5408 2647 5472
rect 2711 5408 2727 5472
rect 2791 5408 2807 5472
rect 2871 5408 2887 5472
rect 2951 5408 2959 5472
rect 2639 4384 2959 5408
rect 2639 4320 2647 4384
rect 2711 4320 2727 4384
rect 2791 4320 2807 4384
rect 2871 4320 2887 4384
rect 2951 4320 2959 4384
rect 2639 3974 2959 4320
rect 2639 3738 2681 3974
rect 2917 3738 2959 3974
rect 2639 3296 2959 3738
rect 2639 3232 2647 3296
rect 2711 3232 2727 3296
rect 2791 3232 2807 3296
rect 2871 3232 2887 3296
rect 2951 3232 2959 3296
rect 2639 2208 2959 3232
rect 2639 2144 2647 2208
rect 2711 2144 2727 2208
rect 2791 2144 2807 2208
rect 2871 2144 2887 2208
rect 2951 2144 2959 2208
rect 2639 2128 2959 2144
rect 4049 10368 4369 10384
rect 4049 10304 4057 10368
rect 4121 10304 4137 10368
rect 4201 10304 4217 10368
rect 4281 10304 4297 10368
rect 4361 10304 4369 10368
rect 4049 9434 4369 10304
rect 4049 9280 4091 9434
rect 4327 9280 4369 9434
rect 4049 9216 4057 9280
rect 4361 9216 4369 9280
rect 4049 9198 4091 9216
rect 4327 9198 4369 9216
rect 4049 8192 4369 9198
rect 4049 8128 4057 8192
rect 4121 8128 4137 8192
rect 4201 8128 4217 8192
rect 4281 8128 4297 8192
rect 4361 8128 4369 8192
rect 4049 7394 4369 8128
rect 4049 7158 4091 7394
rect 4327 7158 4369 7394
rect 4049 7104 4369 7158
rect 4049 7040 4057 7104
rect 4121 7040 4137 7104
rect 4201 7040 4217 7104
rect 4281 7040 4297 7104
rect 4361 7040 4369 7104
rect 4049 6016 4369 7040
rect 4049 5952 4057 6016
rect 4121 5952 4137 6016
rect 4201 5952 4217 6016
rect 4281 5952 4297 6016
rect 4361 5952 4369 6016
rect 4049 5354 4369 5952
rect 4049 5118 4091 5354
rect 4327 5118 4369 5354
rect 4049 4928 4369 5118
rect 4049 4864 4057 4928
rect 4121 4864 4137 4928
rect 4201 4864 4217 4928
rect 4281 4864 4297 4928
rect 4361 4864 4369 4928
rect 4049 3840 4369 4864
rect 4049 3776 4057 3840
rect 4121 3776 4137 3840
rect 4201 3776 4217 3840
rect 4281 3776 4297 3840
rect 4361 3776 4369 3840
rect 4049 3314 4369 3776
rect 4049 3078 4091 3314
rect 4327 3078 4369 3314
rect 4049 2752 4369 3078
rect 4049 2688 4057 2752
rect 4121 2688 4137 2752
rect 4201 2688 4217 2752
rect 4281 2688 4297 2752
rect 4361 2688 4369 2752
rect 4049 2128 4369 2688
rect 4709 10094 5029 10384
rect 4709 9858 4751 10094
rect 4987 9858 5029 10094
rect 4709 9824 5029 9858
rect 4709 9760 4717 9824
rect 4781 9760 4797 9824
rect 4861 9760 4877 9824
rect 4941 9760 4957 9824
rect 5021 9760 5029 9824
rect 4709 8736 5029 9760
rect 4709 8672 4717 8736
rect 4781 8672 4797 8736
rect 4861 8672 4877 8736
rect 4941 8672 4957 8736
rect 5021 8672 5029 8736
rect 4709 8054 5029 8672
rect 4709 7818 4751 8054
rect 4987 7818 5029 8054
rect 4709 7648 5029 7818
rect 4709 7584 4717 7648
rect 4781 7584 4797 7648
rect 4861 7584 4877 7648
rect 4941 7584 4957 7648
rect 5021 7584 5029 7648
rect 4709 6560 5029 7584
rect 4709 6496 4717 6560
rect 4781 6496 4797 6560
rect 4861 6496 4877 6560
rect 4941 6496 4957 6560
rect 5021 6496 5029 6560
rect 4709 6014 5029 6496
rect 4709 5778 4751 6014
rect 4987 5778 5029 6014
rect 4709 5472 5029 5778
rect 4709 5408 4717 5472
rect 4781 5408 4797 5472
rect 4861 5408 4877 5472
rect 4941 5408 4957 5472
rect 5021 5408 5029 5472
rect 4709 4384 5029 5408
rect 4709 4320 4717 4384
rect 4781 4320 4797 4384
rect 4861 4320 4877 4384
rect 4941 4320 4957 4384
rect 5021 4320 5029 4384
rect 4709 3974 5029 4320
rect 4709 3738 4751 3974
rect 4987 3738 5029 3974
rect 4709 3296 5029 3738
rect 4709 3232 4717 3296
rect 4781 3232 4797 3296
rect 4861 3232 4877 3296
rect 4941 3232 4957 3296
rect 5021 3232 5029 3296
rect 4709 2208 5029 3232
rect 4709 2144 4717 2208
rect 4781 2144 4797 2208
rect 4861 2144 4877 2208
rect 4941 2144 4957 2208
rect 5021 2144 5029 2208
rect 4709 2128 5029 2144
rect 6119 10368 6439 10384
rect 6119 10304 6127 10368
rect 6191 10304 6207 10368
rect 6271 10304 6287 10368
rect 6351 10304 6367 10368
rect 6431 10304 6439 10368
rect 6119 9434 6439 10304
rect 6119 9280 6161 9434
rect 6397 9280 6439 9434
rect 6119 9216 6127 9280
rect 6431 9216 6439 9280
rect 6119 9198 6161 9216
rect 6397 9198 6439 9216
rect 6119 8192 6439 9198
rect 6119 8128 6127 8192
rect 6191 8128 6207 8192
rect 6271 8128 6287 8192
rect 6351 8128 6367 8192
rect 6431 8128 6439 8192
rect 6119 7394 6439 8128
rect 6119 7158 6161 7394
rect 6397 7158 6439 7394
rect 6119 7104 6439 7158
rect 6119 7040 6127 7104
rect 6191 7040 6207 7104
rect 6271 7040 6287 7104
rect 6351 7040 6367 7104
rect 6431 7040 6439 7104
rect 6119 6016 6439 7040
rect 6119 5952 6127 6016
rect 6191 5952 6207 6016
rect 6271 5952 6287 6016
rect 6351 5952 6367 6016
rect 6431 5952 6439 6016
rect 6119 5354 6439 5952
rect 6119 5118 6161 5354
rect 6397 5118 6439 5354
rect 6119 4928 6439 5118
rect 6119 4864 6127 4928
rect 6191 4864 6207 4928
rect 6271 4864 6287 4928
rect 6351 4864 6367 4928
rect 6431 4864 6439 4928
rect 6119 3840 6439 4864
rect 6119 3776 6127 3840
rect 6191 3776 6207 3840
rect 6271 3776 6287 3840
rect 6351 3776 6367 3840
rect 6431 3776 6439 3840
rect 6119 3314 6439 3776
rect 6119 3078 6161 3314
rect 6397 3078 6439 3314
rect 6119 2752 6439 3078
rect 6119 2688 6127 2752
rect 6191 2688 6207 2752
rect 6271 2688 6287 2752
rect 6351 2688 6367 2752
rect 6431 2688 6439 2752
rect 6119 2128 6439 2688
rect 6779 10094 7099 10384
rect 6779 9858 6821 10094
rect 7057 9858 7099 10094
rect 6779 9824 7099 9858
rect 6779 9760 6787 9824
rect 6851 9760 6867 9824
rect 6931 9760 6947 9824
rect 7011 9760 7027 9824
rect 7091 9760 7099 9824
rect 6779 8736 7099 9760
rect 6779 8672 6787 8736
rect 6851 8672 6867 8736
rect 6931 8672 6947 8736
rect 7011 8672 7027 8736
rect 7091 8672 7099 8736
rect 6779 8054 7099 8672
rect 6779 7818 6821 8054
rect 7057 7818 7099 8054
rect 6779 7648 7099 7818
rect 6779 7584 6787 7648
rect 6851 7584 6867 7648
rect 6931 7584 6947 7648
rect 7011 7584 7027 7648
rect 7091 7584 7099 7648
rect 6779 6560 7099 7584
rect 6779 6496 6787 6560
rect 6851 6496 6867 6560
rect 6931 6496 6947 6560
rect 7011 6496 7027 6560
rect 7091 6496 7099 6560
rect 6779 6014 7099 6496
rect 6779 5778 6821 6014
rect 7057 5778 7099 6014
rect 6779 5472 7099 5778
rect 6779 5408 6787 5472
rect 6851 5408 6867 5472
rect 6931 5408 6947 5472
rect 7011 5408 7027 5472
rect 7091 5408 7099 5472
rect 6779 4384 7099 5408
rect 6779 4320 6787 4384
rect 6851 4320 6867 4384
rect 6931 4320 6947 4384
rect 7011 4320 7027 4384
rect 7091 4320 7099 4384
rect 6779 3974 7099 4320
rect 6779 3738 6821 3974
rect 7057 3738 7099 3974
rect 6779 3296 7099 3738
rect 6779 3232 6787 3296
rect 6851 3232 6867 3296
rect 6931 3232 6947 3296
rect 7011 3232 7027 3296
rect 7091 3232 7099 3296
rect 6779 2208 7099 3232
rect 6779 2144 6787 2208
rect 6851 2144 6867 2208
rect 6931 2144 6947 2208
rect 7011 2144 7027 2208
rect 7091 2144 7099 2208
rect 6779 2128 7099 2144
rect 8189 10368 8509 10384
rect 8189 10304 8197 10368
rect 8261 10304 8277 10368
rect 8341 10304 8357 10368
rect 8421 10304 8437 10368
rect 8501 10304 8509 10368
rect 8189 9434 8509 10304
rect 8189 9280 8231 9434
rect 8467 9280 8509 9434
rect 8189 9216 8197 9280
rect 8501 9216 8509 9280
rect 8189 9198 8231 9216
rect 8467 9198 8509 9216
rect 8189 8192 8509 9198
rect 8189 8128 8197 8192
rect 8261 8128 8277 8192
rect 8341 8128 8357 8192
rect 8421 8128 8437 8192
rect 8501 8128 8509 8192
rect 8189 7394 8509 8128
rect 8189 7158 8231 7394
rect 8467 7158 8509 7394
rect 8189 7104 8509 7158
rect 8189 7040 8197 7104
rect 8261 7040 8277 7104
rect 8341 7040 8357 7104
rect 8421 7040 8437 7104
rect 8501 7040 8509 7104
rect 8189 6016 8509 7040
rect 8189 5952 8197 6016
rect 8261 5952 8277 6016
rect 8341 5952 8357 6016
rect 8421 5952 8437 6016
rect 8501 5952 8509 6016
rect 8189 5354 8509 5952
rect 8189 5118 8231 5354
rect 8467 5118 8509 5354
rect 8189 4928 8509 5118
rect 8189 4864 8197 4928
rect 8261 4864 8277 4928
rect 8341 4864 8357 4928
rect 8421 4864 8437 4928
rect 8501 4864 8509 4928
rect 8189 3840 8509 4864
rect 8189 3776 8197 3840
rect 8261 3776 8277 3840
rect 8341 3776 8357 3840
rect 8421 3776 8437 3840
rect 8501 3776 8509 3840
rect 8189 3314 8509 3776
rect 8189 3078 8231 3314
rect 8467 3078 8509 3314
rect 8189 2752 8509 3078
rect 8189 2688 8197 2752
rect 8261 2688 8277 2752
rect 8341 2688 8357 2752
rect 8421 2688 8437 2752
rect 8501 2688 8509 2752
rect 8189 2128 8509 2688
rect 8849 10094 9169 10384
rect 8849 9858 8891 10094
rect 9127 9858 9169 10094
rect 8849 9824 9169 9858
rect 8849 9760 8857 9824
rect 8921 9760 8937 9824
rect 9001 9760 9017 9824
rect 9081 9760 9097 9824
rect 9161 9760 9169 9824
rect 8849 8736 9169 9760
rect 8849 8672 8857 8736
rect 8921 8672 8937 8736
rect 9001 8672 9017 8736
rect 9081 8672 9097 8736
rect 9161 8672 9169 8736
rect 8849 8054 9169 8672
rect 8849 7818 8891 8054
rect 9127 7818 9169 8054
rect 8849 7648 9169 7818
rect 8849 7584 8857 7648
rect 8921 7584 8937 7648
rect 9001 7584 9017 7648
rect 9081 7584 9097 7648
rect 9161 7584 9169 7648
rect 8849 6560 9169 7584
rect 8849 6496 8857 6560
rect 8921 6496 8937 6560
rect 9001 6496 9017 6560
rect 9081 6496 9097 6560
rect 9161 6496 9169 6560
rect 8849 6014 9169 6496
rect 8849 5778 8891 6014
rect 9127 5778 9169 6014
rect 8849 5472 9169 5778
rect 8849 5408 8857 5472
rect 8921 5408 8937 5472
rect 9001 5408 9017 5472
rect 9081 5408 9097 5472
rect 9161 5408 9169 5472
rect 8849 4384 9169 5408
rect 8849 4320 8857 4384
rect 8921 4320 8937 4384
rect 9001 4320 9017 4384
rect 9081 4320 9097 4384
rect 9161 4320 9169 4384
rect 8849 3974 9169 4320
rect 8849 3738 8891 3974
rect 9127 3738 9169 3974
rect 8849 3296 9169 3738
rect 8849 3232 8857 3296
rect 8921 3232 8937 3296
rect 9001 3232 9017 3296
rect 9081 3232 9097 3296
rect 9161 3232 9169 3296
rect 8849 2208 9169 3232
rect 8849 2144 8857 2208
rect 8921 2144 8937 2208
rect 9001 2144 9017 2208
rect 9081 2144 9097 2208
rect 9161 2144 9169 2208
rect 8849 2128 9169 2144
<< via4 >>
rect 2021 9280 2257 9434
rect 2021 9216 2051 9280
rect 2051 9216 2067 9280
rect 2067 9216 2131 9280
rect 2131 9216 2147 9280
rect 2147 9216 2211 9280
rect 2211 9216 2227 9280
rect 2227 9216 2257 9280
rect 2021 9198 2257 9216
rect 2021 7158 2257 7394
rect 2021 5118 2257 5354
rect 2021 3078 2257 3314
rect 2681 9858 2917 10094
rect 2681 7818 2917 8054
rect 2681 5778 2917 6014
rect 2681 3738 2917 3974
rect 4091 9280 4327 9434
rect 4091 9216 4121 9280
rect 4121 9216 4137 9280
rect 4137 9216 4201 9280
rect 4201 9216 4217 9280
rect 4217 9216 4281 9280
rect 4281 9216 4297 9280
rect 4297 9216 4327 9280
rect 4091 9198 4327 9216
rect 4091 7158 4327 7394
rect 4091 5118 4327 5354
rect 4091 3078 4327 3314
rect 4751 9858 4987 10094
rect 4751 7818 4987 8054
rect 4751 5778 4987 6014
rect 4751 3738 4987 3974
rect 6161 9280 6397 9434
rect 6161 9216 6191 9280
rect 6191 9216 6207 9280
rect 6207 9216 6271 9280
rect 6271 9216 6287 9280
rect 6287 9216 6351 9280
rect 6351 9216 6367 9280
rect 6367 9216 6397 9280
rect 6161 9198 6397 9216
rect 6161 7158 6397 7394
rect 6161 5118 6397 5354
rect 6161 3078 6397 3314
rect 6821 9858 7057 10094
rect 6821 7818 7057 8054
rect 6821 5778 7057 6014
rect 6821 3738 7057 3974
rect 8231 9280 8467 9434
rect 8231 9216 8261 9280
rect 8261 9216 8277 9280
rect 8277 9216 8341 9280
rect 8341 9216 8357 9280
rect 8357 9216 8421 9280
rect 8421 9216 8437 9280
rect 8437 9216 8467 9280
rect 8231 9198 8467 9216
rect 8231 7158 8467 7394
rect 8231 5118 8467 5354
rect 8231 3078 8467 3314
rect 8891 9858 9127 10094
rect 8891 7818 9127 8054
rect 8891 5778 9127 6014
rect 8891 3738 9127 3974
<< metal5 >>
rect 1056 10094 9432 10136
rect 1056 9858 2681 10094
rect 2917 9858 4751 10094
rect 4987 9858 6821 10094
rect 7057 9858 8891 10094
rect 9127 9858 9432 10094
rect 1056 9816 9432 9858
rect 1056 9434 9432 9476
rect 1056 9198 2021 9434
rect 2257 9198 4091 9434
rect 4327 9198 6161 9434
rect 6397 9198 8231 9434
rect 8467 9198 9432 9434
rect 1056 9156 9432 9198
rect 1056 8054 9432 8096
rect 1056 7818 2681 8054
rect 2917 7818 4751 8054
rect 4987 7818 6821 8054
rect 7057 7818 8891 8054
rect 9127 7818 9432 8054
rect 1056 7776 9432 7818
rect 1056 7394 9432 7436
rect 1056 7158 2021 7394
rect 2257 7158 4091 7394
rect 4327 7158 6161 7394
rect 6397 7158 8231 7394
rect 8467 7158 9432 7394
rect 1056 7116 9432 7158
rect 1056 6014 9432 6056
rect 1056 5778 2681 6014
rect 2917 5778 4751 6014
rect 4987 5778 6821 6014
rect 7057 5778 8891 6014
rect 9127 5778 9432 6014
rect 1056 5736 9432 5778
rect 1056 5354 9432 5396
rect 1056 5118 2021 5354
rect 2257 5118 4091 5354
rect 4327 5118 6161 5354
rect 6397 5118 8231 5354
rect 8467 5118 9432 5354
rect 1056 5076 9432 5118
rect 1056 3974 9432 4016
rect 1056 3738 2681 3974
rect 2917 3738 4751 3974
rect 4987 3738 6821 3974
rect 7057 3738 8891 3974
rect 9127 3738 9432 3974
rect 1056 3696 9432 3738
rect 1056 3314 9432 3356
rect 1056 3078 2021 3314
rect 2257 3078 4091 3314
rect 4327 3078 6161 3314
rect 6397 3078 8231 3314
rect 8467 3078 9432 3314
rect 1056 3036 9432 3078
use sky130_fd_sc_hd__a21oi_1  _084_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 8096 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__or2b_1  _085_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 7728 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _086_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 7912 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _087_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 9016 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _088_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 8924 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  _089_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 7912 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_1  _090_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 7728 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _091_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 6256 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__a21bo_1  _092_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 6256 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__nand3b_1  _093_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 6992 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _094_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 8004 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _095_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 6716 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _096_
timestamp 1723858470
transform 1 0 7820 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _097_
timestamp 1723858470
transform -1 0 8556 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _098_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 7728 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _099_
timestamp 1723858470
transform 1 0 7636 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_2  _100_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 6348 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__or3b_1  _101_
timestamp 1723858470
transform -1 0 7728 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _102_
timestamp 1723858470
transform 1 0 7268 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _103_
timestamp 1723858470
transform -1 0 6992 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _104_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 7636 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _105_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 8280 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _106_
timestamp 1723858470
transform -1 0 8832 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _107_
timestamp 1723858470
transform 1 0 7268 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _108_
timestamp 1723858470
transform 1 0 2760 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_2  _109_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 2484 0 1 7616
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_1  _110_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 4416 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _111_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 6072 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _112_
timestamp 1723858470
transform -1 0 5612 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _113_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 5428 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _114_
timestamp 1723858470
transform -1 0 5888 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _115_
timestamp 1723858470
transform 1 0 5520 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a311o_1  _116_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 4784 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _117_
timestamp 1723858470
transform 1 0 1932 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _118_
timestamp 1723858470
transform 1 0 1656 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _119_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 4508 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _120_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 3772 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _121_
timestamp 1723858470
transform -1 0 4416 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _122_
timestamp 1723858470
transform 1 0 5060 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _123_
timestamp 1723858470
transform 1 0 4416 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _124_
timestamp 1723858470
transform 1 0 3588 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _125_
timestamp 1723858470
transform -1 0 2668 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _126_
timestamp 1723858470
transform -1 0 2944 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a311o_1  _127_
timestamp 1723858470
transform -1 0 3404 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _128_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 3956 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__o41a_1  _129_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 2392 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__xor2_1  _130_
timestamp 1723858470
transform 1 0 1472 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _131_
timestamp 1723858470
transform 1 0 2300 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__o211ai_2  _132_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 3772 0 1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__o21a_1  _133_
timestamp 1723858470
transform 1 0 3864 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _134_
timestamp 1723858470
transform -1 0 3864 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _135_
timestamp 1723858470
transform -1 0 1748 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _136_
timestamp 1723858470
transform 1 0 1748 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _137_
timestamp 1723858470
transform -1 0 2300 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _138_
timestamp 1723858470
transform -1 0 4508 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _139_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 3496 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _140_
timestamp 1723858470
transform -1 0 2668 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _141_
timestamp 1723858470
transform 1 0 2576 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _142_
timestamp 1723858470
transform 1 0 3128 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _143_
timestamp 1723858470
transform 1 0 3220 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _144_
timestamp 1723858470
transform -1 0 4140 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _145_
timestamp 1723858470
transform 1 0 2484 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _146_
timestamp 1723858470
transform 1 0 2668 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _147_
timestamp 1723858470
transform -1 0 4048 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _148_
timestamp 1723858470
transform -1 0 3128 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _149_
timestamp 1723858470
transform 1 0 3128 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _150_
timestamp 1723858470
transform 1 0 1564 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _151_
timestamp 1723858470
transform -1 0 2576 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _152_
timestamp 1723858470
transform 1 0 1748 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _153_
timestamp 1723858470
transform 1 0 1656 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _154_
timestamp 1723858470
transform 1 0 4324 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _155_
timestamp 1723858470
transform 1 0 4048 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _156_
timestamp 1723858470
transform -1 0 5980 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _157_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 5152 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _158_
timestamp 1723858470
transform 1 0 4048 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _159_
timestamp 1723858470
transform -1 0 5152 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _160_
timestamp 1723858470
transform 1 0 4416 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _161_
timestamp 1723858470
transform -1 0 5796 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _162_
timestamp 1723858470
transform -1 0 5980 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _163_
timestamp 1723858470
transform 1 0 5060 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _164_
timestamp 1723858470
transform 1 0 4784 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _165_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 6440 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _166_
timestamp 1723858470
transform -1 0 5796 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__o31a_1  _167_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 5336 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _168_
timestamp 1723858470
transform -1 0 8004 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _169_
timestamp 1723858470
transform 1 0 6624 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _170_
timestamp 1723858470
transform 1 0 6992 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _171_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 7176 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _172_
timestamp 1723858470
transform 1 0 8004 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _173_
timestamp 1723858470
transform 1 0 7360 0 1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _174_
timestamp 1723858470
transform -1 0 7912 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _175_
timestamp 1723858470
transform -1 0 8096 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_7 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 1748 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_33 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 4140 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_45 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 5244 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_55
timestamp 1723858470
transform 1 0 6164 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_57
timestamp 1723858470
transform 1 0 6348 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_65 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 7084 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_79
timestamp 1723858470
transform 1 0 8372 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_85
timestamp 1723858470
transform 1 0 8924 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_3
timestamp 1723858470
transform 1 0 1380 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_29
timestamp 1723858470
transform 1 0 3772 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_53
timestamp 1723858470
transform 1 0 5980 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_57
timestamp 1723858470
transform 1 0 6348 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_77
timestamp 1723858470
transform 1 0 8188 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_14 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 2392 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1723858470
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_29
timestamp 1723858470
transform 1 0 3772 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_39 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 4692 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_50
timestamp 1723858470
transform 1 0 5704 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_62
timestamp 1723858470
transform 1 0 6808 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_75
timestamp 1723858470
transform 1 0 8004 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_79
timestamp 1723858470
transform 1 0 8372 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_83
timestamp 1723858470
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_85
timestamp 1723858470
transform 1 0 8924 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_3
timestamp 1723858470
transform 1 0 1380 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_12
timestamp 1723858470
transform 1 0 2208 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_18
timestamp 1723858470
transform 1 0 2760 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_33
timestamp 1723858470
transform 1 0 4140 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_45
timestamp 1723858470
transform 1 0 5244 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_53
timestamp 1723858470
transform 1 0 5980 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_57
timestamp 1723858470
transform 1 0 6348 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_63
timestamp 1723858470
transform 1 0 6900 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_68
timestamp 1723858470
transform 1 0 7360 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_80
timestamp 1723858470
transform 1 0 8464 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_86
timestamp 1723858470
transform 1 0 9016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_7
timestamp 1723858470
transform 1 0 1748 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_18
timestamp 1723858470
transform 1 0 2760 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_26
timestamp 1723858470
transform 1 0 3496 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_35
timestamp 1723858470
transform 1 0 4324 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_39
timestamp 1723858470
transform 1 0 4692 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_53
timestamp 1723858470
transform 1 0 5980 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_57
timestamp 1723858470
transform 1 0 6348 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_64
timestamp 1723858470
transform 1 0 6992 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_71
timestamp 1723858470
transform 1 0 7636 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_79
timestamp 1723858470
transform 1 0 8372 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_83
timestamp 1723858470
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_85
timestamp 1723858470
transform 1 0 8924 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_14
timestamp 1723858470
transform 1 0 2392 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_22
timestamp 1723858470
transform 1 0 3128 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_34
timestamp 1723858470
transform 1 0 4232 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_51
timestamp 1723858470
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_55
timestamp 1723858470
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_57
timestamp 1723858470
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_76
timestamp 1723858470
transform 1 0 8096 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_3
timestamp 1723858470
transform 1 0 1380 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_20
timestamp 1723858470
transform 1 0 2944 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_29
timestamp 1723858470
transform 1 0 3772 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_37
timestamp 1723858470
transform 1 0 4508 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_44
timestamp 1723858470
transform 1 0 5152 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_56
timestamp 1723858470
transform 1 0 6256 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_64
timestamp 1723858470
transform 1 0 6992 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_78
timestamp 1723858470
transform 1 0 8280 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_85
timestamp 1723858470
transform 1 0 8924 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_3
timestamp 1723858470
transform 1 0 1380 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_17
timestamp 1723858470
transform 1 0 2668 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_44
timestamp 1723858470
transform 1 0 5152 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_72
timestamp 1723858470
transform 1 0 7728 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_86
timestamp 1723858470
transform 1 0 9016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_3
timestamp 1723858470
transform 1 0 1380 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_11
timestamp 1723858470
transform 1 0 2116 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_23
timestamp 1723858470
transform 1 0 3220 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 1723858470
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_39
timestamp 1723858470
transform 1 0 4692 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_51
timestamp 1723858470
transform 1 0 5796 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_63
timestamp 1723858470
transform 1 0 6900 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_80
timestamp 1723858470
transform 1 0 8464 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_85
timestamp 1723858470
transform 1 0 8924 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_9
timestamp 1723858470
transform 1 0 1932 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_13
timestamp 1723858470
transform 1 0 2300 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_23
timestamp 1723858470
transform 1 0 3220 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_35
timestamp 1723858470
transform 1 0 4324 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_43
timestamp 1723858470
transform 1 0 5060 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_49
timestamp 1723858470
transform 1 0 5612 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_55
timestamp 1723858470
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_57
timestamp 1723858470
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_69
timestamp 1723858470
transform 1 0 7452 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_77
timestamp 1723858470
transform 1 0 8188 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_85
timestamp 1723858470
transform 1 0 8924 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_3
timestamp 1723858470
transform 1 0 1380 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_29
timestamp 1723858470
transform 1 0 3772 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_35
timestamp 1723858470
transform 1 0 4324 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_54
timestamp 1723858470
transform 1 0 6072 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_81
timestamp 1723858470
transform 1 0 8556 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_85
timestamp 1723858470
transform 1 0 8924 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_3
timestamp 1723858470
transform 1 0 1380 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_13
timestamp 1723858470
transform 1 0 2300 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_17
timestamp 1723858470
transform 1 0 2668 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_24
timestamp 1723858470
transform 1 0 3312 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_30
timestamp 1723858470
transform 1 0 3864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_38
timestamp 1723858470
transform 1 0 4600 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_47
timestamp 1723858470
transform 1 0 5428 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_55
timestamp 1723858470
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_57
timestamp 1723858470
transform 1 0 6348 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_79
timestamp 1723858470
transform 1 0 8372 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_20
timestamp 1723858470
transform 1 0 2944 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_37
timestamp 1723858470
transform 1 0 4508 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_45
timestamp 1723858470
transform 1 0 5244 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_52
timestamp 1723858470
transform 1 0 5888 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_64
timestamp 1723858470
transform 1 0 6992 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_79
timestamp 1723858470
transform 1 0 8372 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_85
timestamp 1723858470
transform 1 0 8924 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_25
timestamp 1723858470
transform 1 0 3404 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_55
timestamp 1723858470
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_57
timestamp 1723858470
transform 1 0 6348 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_84
timestamp 1723858470
transform 1 0 8832 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_7
timestamp 1723858470
transform 1 0 1748 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_23
timestamp 1723858470
transform 1 0 3220 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_27
timestamp 1723858470
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_29
timestamp 1723858470
transform 1 0 3772 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_37
timestamp 1723858470
transform 1 0 4508 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_44
timestamp 1723858470
transform 1 0 5152 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_57
timestamp 1723858470
transform 1 0 6348 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_65
timestamp 1723858470
transform 1 0 7084 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_77
timestamp 1723858470
transform 1 0 8188 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_85
timestamp 1723858470
transform 1 0 8924 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  input1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 7912 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 9108 0 -1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 5796 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input4
timestamp 1723858470
transform 1 0 1380 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input5
timestamp 1723858470
transform 1 0 1380 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input6
timestamp 1723858470
transform 1 0 1380 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input7
timestamp 1723858470
transform -1 0 7820 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input8
timestamp 1723858470
transform -1 0 8740 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input9
timestamp 1723858470
transform 1 0 2300 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input10
timestamp 1723858470
transform -1 0 8188 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input11
timestamp 1723858470
transform -1 0 8832 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input12
timestamp 1723858470
transform 1 0 1380 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input13
timestamp 1723858470
transform 1 0 1380 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input14
timestamp 1723858470
transform -1 0 8832 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input15
timestamp 1723858470
transform 1 0 1380 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input16
timestamp 1723858470
transform 1 0 2668 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input17
timestamp 1723858470
transform 1 0 2852 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input18
timestamp 1723858470
transform -1 0 9108 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input19
timestamp 1723858470
transform 1 0 3772 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output20 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 8556 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output21
timestamp 1723858470
transform -1 0 8832 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output22
timestamp 1723858470
transform -1 0 5152 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output23
timestamp 1723858470
transform 1 0 6532 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output24
timestamp 1723858470
transform 1 0 6532 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output25
timestamp 1723858470
transform -1 0 1932 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output26
timestamp 1723858470
transform -1 0 2852 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output27
timestamp 1723858470
transform 1 0 8464 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1723858470
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1723858470
transform -1 0 9384 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1723858470
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1723858470
transform -1 0 9384 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1723858470
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1723858470
transform -1 0 9384 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1723858470
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1723858470
transform -1 0 9384 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1723858470
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1723858470
transform -1 0 9384 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1723858470
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1723858470
transform -1 0 9384 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1723858470
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1723858470
transform -1 0 9384 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1723858470
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1723858470
transform -1 0 9384 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1723858470
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1723858470
transform -1 0 9384 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1723858470
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1723858470
transform -1 0 9384 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1723858470
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1723858470
transform -1 0 9384 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1723858470
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1723858470
transform -1 0 9384 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1723858470
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1723858470
transform -1 0 9384 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1723858470
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1723858470
transform -1 0 9384 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1723858470
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1723858470
transform -1 0 9384 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_30 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_31
timestamp 1723858470
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_32
timestamp 1723858470
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_33
timestamp 1723858470
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_34
timestamp 1723858470
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_35
timestamp 1723858470
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_36
timestamp 1723858470
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_37
timestamp 1723858470
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_38
timestamp 1723858470
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_39
timestamp 1723858470
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_40
timestamp 1723858470
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_41
timestamp 1723858470
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_42
timestamp 1723858470
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_43
timestamp 1723858470
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_44
timestamp 1723858470
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_45
timestamp 1723858470
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_46
timestamp 1723858470
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_47
timestamp 1723858470
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_48
timestamp 1723858470
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_49
timestamp 1723858470
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_50
timestamp 1723858470
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_51
timestamp 1723858470
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_52
timestamp 1723858470
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_53
timestamp 1723858470
transform 1 0 6256 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_54
timestamp 1723858470
transform 1 0 8832 0 1 9792
box -38 -48 130 592
<< labels >>
flabel metal4 s 2639 2128 2959 10384 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 4709 2128 5029 10384 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 6779 2128 7099 10384 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 8849 2128 9169 10384 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 3696 9432 4016 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 5736 9432 6056 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 7776 9432 8096 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 9816 9432 10136 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 1979 2128 2299 10384 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 4049 2128 4369 10384 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 6119 2128 6439 10384 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 8189 2128 8509 10384 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 3036 9432 3356 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 5076 9432 5396 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 7116 9432 7436 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 9156 9432 9476 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal3 s 9767 688 10567 808 0 FreeSans 480 0 0 0 a[0]
port 2 nsew signal input
flabel metal3 s 9767 4768 10567 4888 0 FreeSans 480 0 0 0 a[1]
port 3 nsew signal input
flabel metal2 s 5170 0 5226 800 0 FreeSans 224 90 0 0 a[2]
port 4 nsew signal input
flabel metal3 s 0 8848 800 8968 0 FreeSans 480 0 0 0 a[3]
port 5 nsew signal input
flabel metal3 s 0 3408 800 3528 0 FreeSans 480 0 0 0 a[4]
port 6 nsew signal input
flabel metal3 s 0 10208 800 10328 0 FreeSans 480 0 0 0 a[5]
port 7 nsew signal input
flabel metal2 s 9678 11911 9734 12711 0 FreeSans 224 90 0 0 a[6]
port 8 nsew signal input
flabel metal2 s 8390 0 8446 800 0 FreeSans 224 90 0 0 a[7]
port 9 nsew signal input
flabel metal3 s 0 1368 800 1488 0 FreeSans 480 0 0 0 b[0]
port 10 nsew signal input
flabel metal2 s 7746 11911 7802 12711 0 FreeSans 224 90 0 0 b[1]
port 11 nsew signal input
flabel metal3 s 9767 11568 10567 11688 0 FreeSans 480 0 0 0 b[2]
port 12 nsew signal input
flabel metal3 s 0 4768 800 4888 0 FreeSans 480 0 0 0 b[3]
port 13 nsew signal input
flabel metal2 s 1306 11911 1362 12711 0 FreeSans 224 90 0 0 b[4]
port 14 nsew signal input
flabel metal2 s 10322 0 10378 800 0 FreeSans 224 90 0 0 b[5]
port 15 nsew signal input
flabel metal2 s 18 0 74 800 0 FreeSans 224 90 0 0 b[6]
port 16 nsew signal input
flabel metal2 s 1306 0 1362 800 0 FreeSans 224 90 0 0 b[7]
port 17 nsew signal input
flabel metal2 s 2594 11911 2650 12711 0 FreeSans 224 90 0 0 op[0]
port 18 nsew signal input
flabel metal3 s 9767 2728 10567 2848 0 FreeSans 480 0 0 0 op[1]
port 19 nsew signal input
flabel metal2 s 3238 0 3294 800 0 FreeSans 224 90 0 0 op[2]
port 20 nsew signal input
flabel metal3 s 9767 8168 10567 8288 0 FreeSans 480 0 0 0 result[0]
port 21 nsew signal tristate
flabel metal3 s 9767 10208 10567 10328 0 FreeSans 480 0 0 0 result[1]
port 22 nsew signal tristate
flabel metal2 s 4526 11911 4582 12711 0 FreeSans 224 90 0 0 result[2]
port 23 nsew signal tristate
flabel metal2 s 6458 11911 6514 12711 0 FreeSans 224 90 0 0 result[3]
port 24 nsew signal tristate
flabel metal2 s 6458 0 6514 800 0 FreeSans 224 90 0 0 result[4]
port 25 nsew signal tristate
flabel metal3 s 0 6808 800 6928 0 FreeSans 480 0 0 0 result[5]
port 26 nsew signal tristate
flabel metal3 s 0 12248 800 12368 0 FreeSans 480 0 0 0 result[6]
port 27 nsew signal tristate
flabel metal3 s 9767 6128 10567 6248 0 FreeSans 480 0 0 0 result[7]
port 28 nsew signal tristate
rlabel metal1 5244 9792 5244 9792 0 VGND
rlabel metal1 5244 10336 5244 10336 0 VPWR
rlabel metal1 5290 5168 5290 5168 0 _000_
rlabel metal1 5474 5236 5474 5236 0 _001_
rlabel metal2 5382 4862 5382 4862 0 _002_
rlabel metal2 4554 5338 4554 5338 0 _003_
rlabel metal1 5290 4624 5290 4624 0 _004_
rlabel metal1 5704 2618 5704 2618 0 _005_
rlabel metal1 5750 3162 5750 3162 0 _006_
rlabel metal2 5106 4148 5106 4148 0 _007_
rlabel metal1 7130 4658 7130 4658 0 _008_
rlabel metal2 7222 4896 7222 4896 0 _009_
rlabel metal1 6854 3060 6854 3060 0 _010_
rlabel metal1 7176 2958 7176 2958 0 _011_
rlabel metal2 7314 3604 7314 3604 0 _012_
rlabel metal1 7498 3978 7498 3978 0 _013_
rlabel metal1 7728 4794 7728 4794 0 _014_
rlabel metal1 7958 2482 7958 2482 0 _015_
rlabel metal1 7498 2618 7498 2618 0 _016_
rlabel metal1 7728 3162 7728 3162 0 _017_
rlabel metal1 8970 6324 8970 6324 0 _018_
rlabel metal1 8096 5882 8096 5882 0 _019_
rlabel metal1 8648 6222 8648 6222 0 _020_
rlabel metal2 8694 6902 8694 6902 0 _021_
rlabel metal1 6808 9690 6808 9690 0 _022_
rlabel metal1 6210 6358 6210 6358 0 _023_
rlabel viali 6766 7854 6766 7854 0 _024_
rlabel metal1 7038 8602 7038 8602 0 _025_
rlabel metal1 7360 8058 7360 8058 0 _026_
rlabel metal2 7590 8160 7590 8160 0 _027_
rlabel metal1 7222 8534 7222 8534 0 _028_
rlabel metal1 8142 8602 8142 8602 0 _029_
rlabel metal1 7774 8432 7774 8432 0 _030_
rlabel metal1 8464 9078 8464 9078 0 _031_
rlabel metal1 5290 3468 5290 3468 0 _032_
rlabel via1 5750 9554 5750 9554 0 _033_
rlabel metal1 7176 5882 7176 5882 0 _034_
rlabel metal1 1564 5270 1564 5270 0 _035_
rlabel metal1 7314 9520 7314 9520 0 _036_
rlabel metal1 7682 9486 7682 9486 0 _037_
rlabel metal1 8464 9486 8464 9486 0 _038_
rlabel metal2 6026 8126 6026 8126 0 _039_
rlabel metal1 2162 7888 2162 7888 0 _040_
rlabel metal1 4094 7922 4094 7922 0 _041_
rlabel metal1 5842 7888 5842 7888 0 _042_
rlabel metal1 4830 6358 4830 6358 0 _043_
rlabel metal1 5336 7514 5336 7514 0 _044_
rlabel metal1 5336 8602 5336 8602 0 _045_
rlabel metal1 5842 9452 5842 9452 0 _046_
rlabel metal1 5520 9554 5520 9554 0 _047_
rlabel metal1 1886 8058 1886 8058 0 _048_
rlabel metal1 4186 8568 4186 8568 0 _049_
rlabel metal1 4554 9146 4554 9146 0 _050_
rlabel metal2 4324 8942 4324 8942 0 _051_
rlabel metal1 3910 9622 3910 9622 0 _052_
rlabel metal1 4830 9350 4830 9350 0 _053_
rlabel metal1 3680 9622 3680 9622 0 _054_
rlabel metal1 2806 9520 2806 9520 0 _055_
rlabel metal1 2622 9044 2622 9044 0 _056_
rlabel metal2 2714 9350 2714 9350 0 _057_
rlabel metal1 4462 6766 4462 6766 0 _058_
rlabel metal1 2116 6902 2116 6902 0 _059_
rlabel metal1 2392 5746 2392 5746 0 _060_
rlabel metal1 3220 6290 3220 6290 0 _061_
rlabel metal1 4186 5644 4186 5644 0 _062_
rlabel metal1 3864 6290 3864 6290 0 _063_
rlabel metal1 4186 5746 4186 5746 0 _064_
rlabel metal1 2070 5168 2070 5168 0 _065_
rlabel metal2 1794 5508 1794 5508 0 _066_
rlabel metal1 2507 5814 2507 5814 0 _067_
rlabel metal1 3404 3026 3404 3026 0 _068_
rlabel metal1 2990 2958 2990 2958 0 _069_
rlabel metal1 3220 3026 3220 3026 0 _070_
rlabel metal1 4048 4046 4048 4046 0 _071_
rlabel metal1 3910 4046 3910 4046 0 _072_
rlabel metal1 3266 4046 3266 4046 0 _073_
rlabel metal2 2898 4998 2898 4998 0 _074_
rlabel metal1 3450 4590 3450 4590 0 _075_
rlabel metal1 3680 4114 3680 4114 0 _076_
rlabel metal1 2070 4012 2070 4012 0 _077_
rlabel metal1 2162 4046 2162 4046 0 _078_
rlabel metal1 2254 2992 2254 2992 0 _079_
rlabel metal1 2392 3162 2392 3162 0 _080_
rlabel metal1 1840 3706 1840 3706 0 _081_
rlabel metal1 4370 3060 4370 3060 0 _082_
rlabel metal1 5658 4590 5658 4590 0 _083_
rlabel metal3 8932 748 8932 748 0 a[0]
rlabel metal2 9062 4981 9062 4981 0 a[1]
rlabel metal2 5198 823 5198 823 0 a[2]
rlabel metal3 820 8908 820 8908 0 a[3]
rlabel metal3 820 3468 820 3468 0 a[4]
rlabel metal3 1119 10268 1119 10268 0 a[5]
rlabel metal1 8694 9962 8694 9962 0 a[6]
rlabel metal2 8418 823 8418 823 0 a[7]
rlabel metal3 958 1428 958 1428 0 b[0]
rlabel metal1 7912 10030 7912 10030 0 b[1]
rlabel metal1 9062 8942 9062 8942 0 b[2]
rlabel metal3 820 4828 820 4828 0 b[3]
rlabel metal1 1426 10030 1426 10030 0 b[4]
rlabel metal2 10350 1554 10350 1554 0 b[5]
rlabel metal2 46 1554 46 1554 0 b[6]
rlabel metal2 1334 1622 1334 1622 0 b[7]
rlabel metal1 8326 6256 8326 6256 0 net1
rlabel metal1 3220 8262 3220 8262 0 net10
rlabel metal1 2530 7786 2530 7786 0 net11
rlabel metal1 1886 8500 1886 8500 0 net12
rlabel metal1 1794 6766 1794 6766 0 net13
rlabel metal1 5106 2992 5106 2992 0 net14
rlabel metal1 4232 2618 4232 2618 0 net15
rlabel metal1 4945 2482 4945 2482 0 net16
rlabel metal1 4876 9894 4876 9894 0 net17
rlabel metal2 8142 3808 8142 3808 0 net18
rlabel metal1 5382 2550 5382 2550 0 net19
rlabel metal1 8050 7786 8050 7786 0 net2
rlabel metal1 8786 7514 8786 7514 0 net20
rlabel metal1 8740 9622 8740 9622 0 net21
rlabel metal1 4968 9690 4968 9690 0 net22
rlabel metal1 3588 9350 3588 9350 0 net23
rlabel metal1 6256 2414 6256 2414 0 net24
rlabel metal2 1748 7140 1748 7140 0 net25
rlabel metal2 2576 4658 2576 4658 0 net26
rlabel metal2 8050 5508 8050 5508 0 net27
rlabel metal2 6026 2689 6026 2689 0 net3
rlabel metal1 2024 8942 2024 8942 0 net4
rlabel metal1 1564 5202 1564 5202 0 net5
rlabel metal1 1656 3162 1656 3162 0 net6
rlabel metal1 6762 4760 6762 4760 0 net7
rlabel metal1 7498 2482 7498 2482 0 net8
rlabel metal1 3358 7378 3358 7378 0 net9
rlabel metal2 2622 11026 2622 11026 0 op[0]
rlabel metal1 9200 3026 9200 3026 0 op[1]
rlabel metal2 3266 1554 3266 1554 0 op[2]
rlabel metal1 9016 8330 9016 8330 0 result[0]
rlabel metal1 9016 9690 9016 9690 0 result[1]
rlabel metal1 4692 10234 4692 10234 0 result[2]
rlabel metal2 6762 11135 6762 11135 0 result[3]
rlabel metal2 6486 959 6486 959 0 result[4]
rlabel metal3 1096 6868 1096 6868 0 result[5]
rlabel metal3 935 12308 935 12308 0 result[6]
rlabel metal2 8694 6035 8694 6035 0 result[7]
<< properties >>
string FIXED_BBOX 0 0 10567 12711
<< end >>
