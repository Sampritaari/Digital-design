magic
tech sky130A
magscale 1 2
timestamp 1755980430
<< obsli1 >>
rect 1104 2159 9384 10353
<< obsm1 >>
rect 14 2048 10382 10384
<< metal2 >>
rect 1306 11911 1362 12711
rect 2594 11911 2650 12711
rect 4526 11911 4582 12711
rect 6458 11911 6514 12711
rect 7746 11911 7802 12711
rect 9678 11911 9734 12711
rect 18 0 74 800
rect 1306 0 1362 800
rect 3238 0 3294 800
rect 5170 0 5226 800
rect 6458 0 6514 800
rect 8390 0 8446 800
rect 10322 0 10378 800
<< obsm2 >>
rect 20 11855 1250 12050
rect 1418 11855 2538 12050
rect 2706 11855 4470 12050
rect 4638 11855 6402 12050
rect 6570 11855 7690 12050
rect 7858 11855 9622 12050
rect 9790 11855 10376 12050
rect 20 856 10376 11855
rect 130 711 1250 856
rect 1418 711 3182 856
rect 3350 711 5114 856
rect 5282 711 6402 856
rect 6570 711 8334 856
rect 8502 711 10266 856
<< metal3 >>
rect 0 12248 800 12368
rect 9767 11568 10567 11688
rect 0 10208 800 10328
rect 9767 10208 10567 10328
rect 0 8848 800 8968
rect 9767 8168 10567 8288
rect 0 6808 800 6928
rect 9767 6128 10567 6248
rect 0 4768 800 4888
rect 9767 4768 10567 4888
rect 0 3408 800 3528
rect 9767 2728 10567 2848
rect 0 1368 800 1488
rect 9767 688 10567 808
<< obsm3 >>
rect 880 12168 9767 12338
rect 800 11768 9767 12168
rect 800 11488 9687 11768
rect 800 10408 9767 11488
rect 880 10128 9687 10408
rect 800 9048 9767 10128
rect 880 8768 9767 9048
rect 800 8368 9767 8768
rect 800 8088 9687 8368
rect 800 7008 9767 8088
rect 880 6728 9767 7008
rect 800 6328 9767 6728
rect 800 6048 9687 6328
rect 800 4968 9767 6048
rect 880 4688 9687 4968
rect 800 3608 9767 4688
rect 880 3328 9767 3608
rect 800 2928 9767 3328
rect 800 2648 9687 2928
rect 800 1568 9767 2648
rect 880 1288 9767 1568
rect 800 888 9767 1288
rect 800 715 9687 888
<< metal4 >>
rect 1979 2128 2299 10384
rect 2639 2128 2959 10384
rect 4049 2128 4369 10384
rect 4709 2128 5029 10384
rect 6119 2128 6439 10384
rect 6779 2128 7099 10384
rect 8189 2128 8509 10384
rect 8849 2128 9169 10384
<< metal5 >>
rect 1056 9816 9432 10136
rect 1056 9156 9432 9476
rect 1056 7776 9432 8096
rect 1056 7116 9432 7436
rect 1056 5736 9432 6056
rect 1056 5076 9432 5396
rect 1056 3696 9432 4016
rect 1056 3036 9432 3356
<< labels >>
rlabel metal4 s 2639 2128 2959 10384 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 4709 2128 5029 10384 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 6779 2128 7099 10384 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 8849 2128 9169 10384 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 3696 9432 4016 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 5736 9432 6056 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 7776 9432 8096 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 9816 9432 10136 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 1979 2128 2299 10384 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 4049 2128 4369 10384 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 6119 2128 6439 10384 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 8189 2128 8509 10384 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 3036 9432 3356 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 5076 9432 5396 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 7116 9432 7436 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 9156 9432 9476 6 VPWR
port 2 nsew power bidirectional
rlabel metal3 s 9767 688 10567 808 6 a[0]
port 3 nsew signal input
rlabel metal3 s 9767 4768 10567 4888 6 a[1]
port 4 nsew signal input
rlabel metal2 s 5170 0 5226 800 6 a[2]
port 5 nsew signal input
rlabel metal3 s 0 8848 800 8968 6 a[3]
port 6 nsew signal input
rlabel metal3 s 0 3408 800 3528 6 a[4]
port 7 nsew signal input
rlabel metal3 s 0 10208 800 10328 6 a[5]
port 8 nsew signal input
rlabel metal2 s 9678 11911 9734 12711 6 a[6]
port 9 nsew signal input
rlabel metal2 s 8390 0 8446 800 6 a[7]
port 10 nsew signal input
rlabel metal3 s 0 1368 800 1488 6 b[0]
port 11 nsew signal input
rlabel metal2 s 7746 11911 7802 12711 6 b[1]
port 12 nsew signal input
rlabel metal3 s 9767 11568 10567 11688 6 b[2]
port 13 nsew signal input
rlabel metal3 s 0 4768 800 4888 6 b[3]
port 14 nsew signal input
rlabel metal2 s 1306 11911 1362 12711 6 b[4]
port 15 nsew signal input
rlabel metal2 s 10322 0 10378 800 6 b[5]
port 16 nsew signal input
rlabel metal2 s 18 0 74 800 6 b[6]
port 17 nsew signal input
rlabel metal2 s 1306 0 1362 800 6 b[7]
port 18 nsew signal input
rlabel metal2 s 2594 11911 2650 12711 6 op[0]
port 19 nsew signal input
rlabel metal3 s 9767 2728 10567 2848 6 op[1]
port 20 nsew signal input
rlabel metal2 s 3238 0 3294 800 6 op[2]
port 21 nsew signal input
rlabel metal3 s 9767 8168 10567 8288 6 result[0]
port 22 nsew signal output
rlabel metal3 s 9767 10208 10567 10328 6 result[1]
port 23 nsew signal output
rlabel metal2 s 4526 11911 4582 12711 6 result[2]
port 24 nsew signal output
rlabel metal2 s 6458 11911 6514 12711 6 result[3]
port 25 nsew signal output
rlabel metal2 s 6458 0 6514 800 6 result[4]
port 26 nsew signal output
rlabel metal3 s 0 6808 800 6928 6 result[5]
port 27 nsew signal output
rlabel metal3 s 0 12248 800 12368 6 result[6]
port 28 nsew signal output
rlabel metal3 s 9767 6128 10567 6248 6 result[7]
port 29 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 10567 12711
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 560380
string GDS_FILE /openlane/designs/alu/runs/RUN_2025.08.23_20.19.57/results/signoff/alu.magic.gds
string GDS_START 223484
<< end >>

