module alu (a,
    b,
    op,
    result);
 input [7:0] a;
 input [7:0] b;
 input [2:0] op;
 output [7:0] result;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;

 sky130_fd_sc_hd__a21oi_2 _084_ (.A1(a[0]),
    .A2(b[0]),
    .B1(op[0]),
    .Y(_018_));
 sky130_fd_sc_hd__or2b_2 _085_ (.A(op[2]),
    .B_N(op[1]),
    .X(_019_));
 sky130_fd_sc_hd__a221o_2 _086_ (.A1(a[0]),
    .A2(b[0]),
    .B1(op[2]),
    .B2(op[0]),
    .C1(op[1]),
    .X(_020_));
 sky130_fd_sc_hd__o21ai_2 _087_ (.A1(_018_),
    .A2(_019_),
    .B1(_020_),
    .Y(_021_));
 sky130_fd_sc_hd__o21a_2 _088_ (.A1(a[0]),
    .A2(b[0]),
    .B1(_021_),
    .X(result[0]));
 sky130_fd_sc_hd__nor2_2 _089_ (.A(op[2]),
    .B(op[1]),
    .Y(_022_));
 sky130_fd_sc_hd__or3b_2 _090_ (.A(op[2]),
    .B(op[1]),
    .C_N(op[0]),
    .X(_023_));
 sky130_fd_sc_hd__buf_1 _091_ (.A(_023_),
    .X(_024_));
 sky130_fd_sc_hd__a21bo_2 _092_ (.A1(b[0]),
    .A2(_024_),
    .B1_N(b[1]),
    .X(_025_));
 sky130_fd_sc_hd__nand3b_2 _093_ (.A_N(b[1]),
    .B(_024_),
    .C(b[0]),
    .Y(_026_));
 sky130_fd_sc_hd__and3_2 _094_ (.A(a[1]),
    .B(_025_),
    .C(_026_),
    .X(_027_));
 sky130_fd_sc_hd__a21o_2 _095_ (.A1(_025_),
    .A2(_026_),
    .B1(a[1]),
    .X(_028_));
 sky130_fd_sc_hd__or2b_2 _096_ (.A(_027_),
    .B_N(_028_),
    .X(_029_));
 sky130_fd_sc_hd__or2b_2 _097_ (.A(a[0]),
    .B_N(b[0]),
    .X(_030_));
 sky130_fd_sc_hd__xnor2_2 _098_ (.A(_029_),
    .B(_030_),
    .Y(_031_));
 sky130_fd_sc_hd__nor2_2 _099_ (.A(op[0]),
    .B(_019_),
    .Y(_032_));
 sky130_fd_sc_hd__and3b_2 _100_ (.A_N(op[2]),
    .B(op[1]),
    .C(op[0]),
    .X(_033_));
 sky130_fd_sc_hd__or3b_2 _101_ (.A(op[1]),
    .B(op[0]),
    .C_N(op[2]),
    .X(_034_));
 sky130_fd_sc_hd__buf_1 _102_ (.A(_034_),
    .X(_035_));
 sky130_fd_sc_hd__a21oi_2 _103_ (.A1(a[1]),
    .A2(b[1]),
    .B1(_035_),
    .Y(_036_));
 sky130_fd_sc_hd__o22a_2 _104_ (.A1(a[1]),
    .A2(b[1]),
    .B1(_033_),
    .B2(_036_),
    .X(_037_));
 sky130_fd_sc_hd__a31o_2 _105_ (.A1(a[1]),
    .A2(b[1]),
    .A3(_032_),
    .B1(_037_),
    .X(_038_));
 sky130_fd_sc_hd__a21o_2 _106_ (.A1(_022_),
    .A2(_031_),
    .B1(_038_),
    .X(result[1]));
 sky130_fd_sc_hd__a21o_2 _107_ (.A1(_028_),
    .A2(_030_),
    .B1(_027_),
    .X(_039_));
 sky130_fd_sc_hd__o21a_2 _108_ (.A1(b[0]),
    .A2(b[1]),
    .B1(_024_),
    .X(_040_));
 sky130_fd_sc_hd__xnor2_2 _109_ (.A(b[2]),
    .B(_040_),
    .Y(_041_));
 sky130_fd_sc_hd__xor2_2 _110_ (.A(a[2]),
    .B(_041_),
    .X(_042_));
 sky130_fd_sc_hd__and2_2 _111_ (.A(_039_),
    .B(_042_),
    .X(_043_));
 sky130_fd_sc_hd__o21ai_2 _112_ (.A1(_039_),
    .A2(_042_),
    .B1(_022_),
    .Y(_044_));
 sky130_fd_sc_hd__nor2_2 _113_ (.A(_043_),
    .B(_044_),
    .Y(_045_));
 sky130_fd_sc_hd__a21oi_2 _114_ (.A1(a[2]),
    .A2(b[2]),
    .B1(_035_),
    .Y(_046_));
 sky130_fd_sc_hd__o22a_2 _115_ (.A1(a[2]),
    .A2(b[2]),
    .B1(_033_),
    .B2(_046_),
    .X(_047_));
 sky130_fd_sc_hd__a311o_2 _116_ (.A1(a[2]),
    .A2(b[2]),
    .A3(_032_),
    .B1(_045_),
    .C1(_047_),
    .X(result[2]));
 sky130_fd_sc_hd__a21o_2 _117_ (.A1(b[2]),
    .A2(_024_),
    .B1(_040_),
    .X(_048_));
 sky130_fd_sc_hd__xnor2_2 _118_ (.A(b[3]),
    .B(_048_),
    .Y(_049_));
 sky130_fd_sc_hd__nand2_2 _119_ (.A(a[3]),
    .B(_049_),
    .Y(_050_));
 sky130_fd_sc_hd__or2_2 _120_ (.A(a[3]),
    .B(_049_),
    .X(_051_));
 sky130_fd_sc_hd__and2_2 _121_ (.A(_050_),
    .B(_051_),
    .X(_052_));
 sky130_fd_sc_hd__a21o_2 _122_ (.A1(a[2]),
    .A2(_041_),
    .B1(_043_),
    .X(_053_));
 sky130_fd_sc_hd__o21ai_2 _123_ (.A1(_052_),
    .A2(_053_),
    .B1(_022_),
    .Y(_054_));
 sky130_fd_sc_hd__a21oi_2 _124_ (.A1(_052_),
    .A2(_053_),
    .B1(_054_),
    .Y(_055_));
 sky130_fd_sc_hd__a21oi_2 _125_ (.A1(a[3]),
    .A2(b[3]),
    .B1(_035_),
    .Y(_056_));
 sky130_fd_sc_hd__o22a_2 _126_ (.A1(a[3]),
    .A2(b[3]),
    .B1(_033_),
    .B2(_056_),
    .X(_057_));
 sky130_fd_sc_hd__a311o_2 _127_ (.A1(a[3]),
    .A2(b[3]),
    .A3(_032_),
    .B1(_055_),
    .C1(_057_),
    .X(result[3]));
 sky130_fd_sc_hd__a22o_2 _128_ (.A1(a[2]),
    .A2(_041_),
    .B1(_049_),
    .B2(a[3]),
    .X(_058_));
 sky130_fd_sc_hd__o41a_2 _129_ (.A1(b[0]),
    .A2(b[1]),
    .A3(b[2]),
    .A4(b[3]),
    .B1(_024_),
    .X(_059_));
 sky130_fd_sc_hd__xor2_2 _130_ (.A(b[4]),
    .B(_059_),
    .X(_060_));
 sky130_fd_sc_hd__xnor2_2 _131_ (.A(a[4]),
    .B(_060_),
    .Y(_061_));
 sky130_fd_sc_hd__o211ai_2 _132_ (.A1(_043_),
    .A2(_058_),
    .B1(_061_),
    .C1(_051_),
    .Y(_062_));
 sky130_fd_sc_hd__o21a_2 _133_ (.A1(_043_),
    .A2(_058_),
    .B1(_051_),
    .X(_063_));
 sky130_fd_sc_hd__or2_2 _134_ (.A(_061_),
    .B(_063_),
    .X(_064_));
 sky130_fd_sc_hd__a21oi_2 _135_ (.A1(a[4]),
    .A2(b[4]),
    .B1(_035_),
    .Y(_065_));
 sky130_fd_sc_hd__o22a_2 _136_ (.A1(a[4]),
    .A2(b[4]),
    .B1(_033_),
    .B2(_065_),
    .X(_066_));
 sky130_fd_sc_hd__a31o_2 _137_ (.A1(a[4]),
    .A2(b[4]),
    .A3(_032_),
    .B1(_066_),
    .X(_067_));
 sky130_fd_sc_hd__a31o_2 _138_ (.A1(_022_),
    .A2(_062_),
    .A3(_064_),
    .B1(_067_),
    .X(result[4]));
 sky130_fd_sc_hd__inv_2 _139_ (.A(a[5]),
    .Y(_068_));
 sky130_fd_sc_hd__a21o_2 _140_ (.A1(b[4]),
    .A2(_024_),
    .B1(_059_),
    .X(_069_));
 sky130_fd_sc_hd__xor2_2 _141_ (.A(b[5]),
    .B(_069_),
    .X(_070_));
 sky130_fd_sc_hd__or2_2 _142_ (.A(_068_),
    .B(_070_),
    .X(_071_));
 sky130_fd_sc_hd__nand2_2 _143_ (.A(_068_),
    .B(_070_),
    .Y(_072_));
 sky130_fd_sc_hd__and2_2 _144_ (.A(_071_),
    .B(_072_),
    .X(_073_));
 sky130_fd_sc_hd__inv_2 _145_ (.A(a[4]),
    .Y(_074_));
 sky130_fd_sc_hd__or2_2 _146_ (.A(_074_),
    .B(_060_),
    .X(_075_));
 sky130_fd_sc_hd__nand2_2 _147_ (.A(_075_),
    .B(_062_),
    .Y(_076_));
 sky130_fd_sc_hd__nand2_2 _148_ (.A(_073_),
    .B(_076_),
    .Y(_077_));
 sky130_fd_sc_hd__o21a_2 _149_ (.A1(_073_),
    .A2(_076_),
    .B1(_022_),
    .X(_078_));
 sky130_fd_sc_hd__a21oi_2 _150_ (.A1(a[5]),
    .A2(b[5]),
    .B1(_035_),
    .Y(_079_));
 sky130_fd_sc_hd__o22a_2 _151_ (.A1(a[5]),
    .A2(b[5]),
    .B1(_033_),
    .B2(_079_),
    .X(_080_));
 sky130_fd_sc_hd__a31o_2 _152_ (.A1(a[5]),
    .A2(b[5]),
    .A3(_032_),
    .B1(_080_),
    .X(_081_));
 sky130_fd_sc_hd__a21o_2 _153_ (.A1(_077_),
    .A2(_078_),
    .B1(_081_),
    .X(result[5]));
 sky130_fd_sc_hd__a21oi_2 _154_ (.A1(b[5]),
    .A2(_024_),
    .B1(_069_),
    .Y(_082_));
 sky130_fd_sc_hd__xnor2_2 _155_ (.A(b[6]),
    .B(_082_),
    .Y(_083_));
 sky130_fd_sc_hd__xnor2_2 _156_ (.A(a[6]),
    .B(_083_),
    .Y(_000_));
 sky130_fd_sc_hd__o211a_2 _157_ (.A1(_043_),
    .A2(_058_),
    .B1(_061_),
    .C1(_051_),
    .X(_001_));
 sky130_fd_sc_hd__nand2_2 _158_ (.A(_075_),
    .B(_071_),
    .Y(_002_));
 sky130_fd_sc_hd__o21ai_2 _159_ (.A1(_001_),
    .A2(_002_),
    .B1(_072_),
    .Y(_003_));
 sky130_fd_sc_hd__xnor2_2 _160_ (.A(_000_),
    .B(_003_),
    .Y(_004_));
 sky130_fd_sc_hd__a21oi_2 _161_ (.A1(a[6]),
    .A2(b[6]),
    .B1(_035_),
    .Y(_005_));
 sky130_fd_sc_hd__o22a_2 _162_ (.A1(a[6]),
    .A2(b[6]),
    .B1(_033_),
    .B2(_005_),
    .X(_006_));
 sky130_fd_sc_hd__a31o_2 _163_ (.A1(a[6]),
    .A2(b[6]),
    .A3(_032_),
    .B1(_006_),
    .X(_007_));
 sky130_fd_sc_hd__a21o_2 _164_ (.A1(_022_),
    .A2(_004_),
    .B1(_007_),
    .X(result[6]));
 sky130_fd_sc_hd__and2b_2 _165_ (.A_N(_083_),
    .B(a[6]),
    .X(_008_));
 sky130_fd_sc_hd__o211a_2 _166_ (.A1(_001_),
    .A2(_002_),
    .B1(_000_),
    .C1(_072_),
    .X(_009_));
 sky130_fd_sc_hd__o31a_2 _167_ (.A1(b[5]),
    .A2(b[6]),
    .A3(_069_),
    .B1(_024_),
    .X(_010_));
 sky130_fd_sc_hd__xor2_2 _168_ (.A(a[7]),
    .B(b[7]),
    .X(_011_));
 sky130_fd_sc_hd__xnor2_2 _169_ (.A(_010_),
    .B(_011_),
    .Y(_012_));
 sky130_fd_sc_hd__o21ai_2 _170_ (.A1(_008_),
    .A2(_009_),
    .B1(_012_),
    .Y(_013_));
 sky130_fd_sc_hd__or3_2 _171_ (.A(_008_),
    .B(_009_),
    .C(_012_),
    .X(_014_));
 sky130_fd_sc_hd__a21oi_2 _172_ (.A1(a[7]),
    .A2(b[7]),
    .B1(_035_),
    .Y(_015_));
 sky130_fd_sc_hd__a31o_2 _173_ (.A1(a[7]),
    .A2(b[7]),
    .A3(_032_),
    .B1(_015_),
    .X(_016_));
 sky130_fd_sc_hd__o22a_2 _174_ (.A1(a[7]),
    .A2(b[7]),
    .B1(_033_),
    .B2(_016_),
    .X(_017_));
 sky130_fd_sc_hd__a31o_2 _175_ (.A1(_022_),
    .A2(_013_),
    .A3(_014_),
    .B1(_017_),
    .X(result[7]));
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_37 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_38 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_39 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_40 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_41 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_42 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_43 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_44 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_45 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_46 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_47 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_48 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_49 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_50 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_51 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_52 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_53 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_54 ();
endmodule
